*
* MAIN CELL: Component pathname : root_element
*
   .MODEL MMI_switch_ideal "label 1"="TE" "control"=1
   .MODEL "Waveguide Crossing" "label 1"="TE" "transmission 1"=0.9954054174 "cross talk 1"=0.0001
   + "transmission 2"=1 "cross talk 2"=0 "reflection 1"=0.001
   + "reflection 2"=0 "label 2"="TM" "orthogonal identifier 1"=1
   + "orthogonal identifier 2"=2
   .MODEL "Straight Waveguide" "excess loss temperature sensitivity 2"=0 "label 1"="TE" "orthogonal identifier 1"=1 
   + "loss 1"=0 "number of taps"=64 "dispersion 1"=0 
   + "effective index temperature sensitivity 2"=0 "effective index 2"=1 length=10u 
   + "group index 2"=1 "orthogonal identifier 2"=2 "nominal temperature"=300 
   + "loss 2"=0 "dispersion 2"=0 frequency=193.1T 
   + "digital filter"=0 "run diagnostic"=0 "window function"="rectangular" 
   + "thermal fill factor"=1 "excess loss temperature sensitivity 1"=0 "label 2"="TM" 
   + "thermal effects"=0 "effective index temperature sensitivity 1"=0 "effective index 1"=1 

.subckt HDBE  N$8961 N$8963 N$8965 N$8967 N$8969 N$8971 N$8973 N$8975 N$8977 N$8979 N$8981 N$8983 N$8985 N$8987 N$8989 N$8991 N$8993 N$8995 N$8997 N$8999 N$9001 N$9003 N$9005 N$9007 N$9009 N$9011 N$9013 N$9015 N$9017 N$9019 N$9021 N$9023 N$9153 N$9155 N$9157 N$9159 N$9161 N$9163 N$9165 N$9167 N$9169 N$9171 N$9173 N$9175 N$9177 N$9179 N$9181 N$9183 N$9185 N$9187 N$9189 N$9191 N$9193 N$9195 N$9197 N$9199 N$9201 N$9203 N$9205 N$9207 N$9209 N$9211 N$9213 N$9215
   S1249 N$8961 N$8962 N$6845 N$4738 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1250 N$8963 N$8964 N$4740 N$4742 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1251 N$8965 N$8966 N$4744 N$4746 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1252 N$8967 N$8968 N$4748 N$4750 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1253 N$8969 N$8970 N$4752 N$4754 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1254 N$8971 N$8972 N$4756 N$4758 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1255 N$8973 N$8974 N$4760 N$4762 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1256 N$8975 N$8976 N$4764 N$4766 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1257 N$8977 N$8978 N$4768 N$4770 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1258 N$8979 N$8980 N$4772 N$4774 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1259 N$8981 N$8982 N$4776 N$4778 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1260 N$8983 N$8984 N$4780 N$4782 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1261 N$8985 N$8986 N$4784 N$4786 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1262 N$8987 N$8988 N$4788 N$4790 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1263 N$8989 N$8990 N$4792 N$4794 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1264 N$8991 N$8992 N$4796 N$4798 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1265 N$8993 N$8994 N$4800 N$4802 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1266 N$8995 N$8996 N$4804 N$4806 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1267 N$8997 N$8998 N$4808 N$4810 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1268 N$8999 N$9000 N$4812 N$4814 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1269 N$9001 N$9002 N$4816 N$4818 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1270 N$9003 N$9004 N$4820 N$4822 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1271 N$9005 N$9006 N$4824 N$4826 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1272 N$9007 N$9008 N$4828 N$4830 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1273 N$9009 N$9010 N$4832 N$4834 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1274 N$9011 N$9012 N$4836 N$4838 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1275 N$9013 N$9014 N$4840 N$4842 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1276 N$9015 N$9016 N$4844 N$4846 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1277 N$9017 N$9018 N$4848 N$4850 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1278 N$9019 N$9020 N$4852 N$4854 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1279 N$9021 N$9022 N$4856 N$4858 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1280 N$9023 N$9024 N$4860 N$6847 MMI_switch_ideal library="Design kits/capstone" sch_x=-126 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1281 N$4737 N$4739 N$6721 N$4862 "Waveguide Crossing" sch_x=-124 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1282 N$4741 N$4743 N$4864 N$4866 "Waveguide Crossing" sch_x=-124 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1283 N$4745 N$4747 N$4868 N$4870 "Waveguide Crossing" sch_x=-124 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1284 N$4749 N$4751 N$4872 N$4874 "Waveguide Crossing" sch_x=-124 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1285 N$4753 N$4755 N$4876 N$4878 "Waveguide Crossing" sch_x=-124 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1286 N$4757 N$4759 N$4880 N$4882 "Waveguide Crossing" sch_x=-124 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1287 N$4761 N$4763 N$4884 N$4886 "Waveguide Crossing" sch_x=-124 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1288 N$4765 N$4767 N$4888 N$4890 "Waveguide Crossing" sch_x=-124 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1289 N$4769 N$4771 N$4892 N$4894 "Waveguide Crossing" sch_x=-124 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1290 N$4773 N$4775 N$4896 N$4898 "Waveguide Crossing" sch_x=-124 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1291 N$4777 N$4779 N$4900 N$4902 "Waveguide Crossing" sch_x=-124 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1292 N$4781 N$4783 N$4904 N$4906 "Waveguide Crossing" sch_x=-124 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1293 N$4785 N$4787 N$4908 N$4910 "Waveguide Crossing" sch_x=-124 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1294 N$4789 N$4791 N$4912 N$4914 "Waveguide Crossing" sch_x=-124 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1295 N$4793 N$4795 N$4916 N$4918 "Waveguide Crossing" sch_x=-124 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1296 N$4797 N$4799 N$4920 N$4922 "Waveguide Crossing" sch_x=-124 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1297 N$4801 N$4803 N$4924 N$4926 "Waveguide Crossing" sch_x=-124 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1298 N$4805 N$4807 N$4928 N$4930 "Waveguide Crossing" sch_x=-124 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1299 N$4809 N$4811 N$4932 N$4934 "Waveguide Crossing" sch_x=-124 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1300 N$4813 N$4815 N$4936 N$4938 "Waveguide Crossing" sch_x=-124 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1301 N$4817 N$4819 N$4940 N$4942 "Waveguide Crossing" sch_x=-124 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1302 N$4821 N$4823 N$4944 N$4946 "Waveguide Crossing" sch_x=-124 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1303 N$4825 N$4827 N$4948 N$4950 "Waveguide Crossing" sch_x=-124 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1304 N$4829 N$4831 N$4952 N$4954 "Waveguide Crossing" sch_x=-124 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1305 N$4833 N$4835 N$4956 N$4958 "Waveguide Crossing" sch_x=-124 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1306 N$4837 N$4839 N$4960 N$4962 "Waveguide Crossing" sch_x=-124 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1307 N$4841 N$4843 N$4964 N$4966 "Waveguide Crossing" sch_x=-124 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1308 N$4845 N$4847 N$4968 N$4970 "Waveguide Crossing" sch_x=-124 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1309 N$4849 N$4851 N$4972 N$4974 "Waveguide Crossing" sch_x=-124 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1310 N$4853 N$4855 N$4976 N$4978 "Waveguide Crossing" sch_x=-124 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1311 N$4857 N$4859 N$4980 N$6843 "Waveguide Crossing" sch_x=-124 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1312 N$4861 N$4863 N$6723 N$4982 "Waveguide Crossing" sch_x=-122 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1313 N$4865 N$4867 N$4984 N$4986 "Waveguide Crossing" sch_x=-122 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1314 N$4869 N$4871 N$4988 N$4990 "Waveguide Crossing" sch_x=-122 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1315 N$4873 N$4875 N$4992 N$4994 "Waveguide Crossing" sch_x=-122 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1316 N$4877 N$4879 N$4996 N$4998 "Waveguide Crossing" sch_x=-122 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1317 N$4881 N$4883 N$5000 N$5002 "Waveguide Crossing" sch_x=-122 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1318 N$4885 N$4887 N$5004 N$5006 "Waveguide Crossing" sch_x=-122 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1319 N$4889 N$4891 N$5008 N$5010 "Waveguide Crossing" sch_x=-122 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1320 N$4893 N$4895 N$5012 N$5014 "Waveguide Crossing" sch_x=-122 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1321 N$4897 N$4899 N$5016 N$5018 "Waveguide Crossing" sch_x=-122 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1322 N$4901 N$4903 N$5020 N$5022 "Waveguide Crossing" sch_x=-122 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1323 N$4905 N$4907 N$5024 N$5026 "Waveguide Crossing" sch_x=-122 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1324 N$4909 N$4911 N$5028 N$5030 "Waveguide Crossing" sch_x=-122 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1325 N$4913 N$4915 N$5032 N$5034 "Waveguide Crossing" sch_x=-122 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1326 N$4917 N$4919 N$5036 N$5038 "Waveguide Crossing" sch_x=-122 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1327 N$4921 N$4923 N$5040 N$5042 "Waveguide Crossing" sch_x=-122 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1328 N$4925 N$4927 N$5044 N$5046 "Waveguide Crossing" sch_x=-122 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1329 N$4929 N$4931 N$5048 N$5050 "Waveguide Crossing" sch_x=-122 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1330 N$4933 N$4935 N$5052 N$5054 "Waveguide Crossing" sch_x=-122 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1331 N$4937 N$4939 N$5056 N$5058 "Waveguide Crossing" sch_x=-122 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1332 N$4941 N$4943 N$5060 N$5062 "Waveguide Crossing" sch_x=-122 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1333 N$4945 N$4947 N$5064 N$5066 "Waveguide Crossing" sch_x=-122 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1334 N$4949 N$4951 N$5068 N$5070 "Waveguide Crossing" sch_x=-122 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1335 N$4953 N$4955 N$5072 N$5074 "Waveguide Crossing" sch_x=-122 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1336 N$4957 N$4959 N$5076 N$5078 "Waveguide Crossing" sch_x=-122 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1337 N$4961 N$4963 N$5080 N$5082 "Waveguide Crossing" sch_x=-122 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1338 N$4965 N$4967 N$5084 N$5086 "Waveguide Crossing" sch_x=-122 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1339 N$4969 N$4971 N$5088 N$5090 "Waveguide Crossing" sch_x=-122 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1340 N$4973 N$4975 N$5092 N$5094 "Waveguide Crossing" sch_x=-122 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1341 N$4977 N$4979 N$5096 N$6841 "Waveguide Crossing" sch_x=-122 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1342 N$4981 N$4983 N$6725 N$5098 "Waveguide Crossing" sch_x=-120 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1343 N$4985 N$4987 N$5100 N$5102 "Waveguide Crossing" sch_x=-120 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1344 N$4989 N$4991 N$5104 N$5106 "Waveguide Crossing" sch_x=-120 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1345 N$4993 N$4995 N$5108 N$5110 "Waveguide Crossing" sch_x=-120 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1346 N$4997 N$4999 N$5112 N$5114 "Waveguide Crossing" sch_x=-120 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1347 N$5001 N$5003 N$5116 N$5118 "Waveguide Crossing" sch_x=-120 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1348 N$5005 N$5007 N$5120 N$5122 "Waveguide Crossing" sch_x=-120 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1349 N$5009 N$5011 N$5124 N$5126 "Waveguide Crossing" sch_x=-120 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1350 N$5013 N$5015 N$5128 N$5130 "Waveguide Crossing" sch_x=-120 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1351 N$5017 N$5019 N$5132 N$5134 "Waveguide Crossing" sch_x=-120 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1352 N$5021 N$5023 N$5136 N$5138 "Waveguide Crossing" sch_x=-120 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1353 N$5025 N$5027 N$5140 N$5142 "Waveguide Crossing" sch_x=-120 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1354 N$5029 N$5031 N$5144 N$5146 "Waveguide Crossing" sch_x=-120 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1355 N$5033 N$5035 N$5148 N$5150 "Waveguide Crossing" sch_x=-120 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1356 N$5037 N$5039 N$5152 N$5154 "Waveguide Crossing" sch_x=-120 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1357 N$5041 N$5043 N$5156 N$5158 "Waveguide Crossing" sch_x=-120 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1358 N$5045 N$5047 N$5160 N$5162 "Waveguide Crossing" sch_x=-120 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1359 N$5049 N$5051 N$5164 N$5166 "Waveguide Crossing" sch_x=-120 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1360 N$5053 N$5055 N$5168 N$5170 "Waveguide Crossing" sch_x=-120 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1361 N$5057 N$5059 N$5172 N$5174 "Waveguide Crossing" sch_x=-120 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1362 N$5061 N$5063 N$5176 N$5178 "Waveguide Crossing" sch_x=-120 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1363 N$5065 N$5067 N$5180 N$5182 "Waveguide Crossing" sch_x=-120 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1364 N$5069 N$5071 N$5184 N$5186 "Waveguide Crossing" sch_x=-120 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1365 N$5073 N$5075 N$5188 N$5190 "Waveguide Crossing" sch_x=-120 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1366 N$5077 N$5079 N$5192 N$5194 "Waveguide Crossing" sch_x=-120 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1367 N$5081 N$5083 N$5196 N$5198 "Waveguide Crossing" sch_x=-120 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1368 N$5085 N$5087 N$5200 N$5202 "Waveguide Crossing" sch_x=-120 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1369 N$5089 N$5091 N$5204 N$5206 "Waveguide Crossing" sch_x=-120 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1370 N$5093 N$5095 N$5208 N$6839 "Waveguide Crossing" sch_x=-120 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1371 N$5097 N$5099 N$6727 N$5210 "Waveguide Crossing" sch_x=-118 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1372 N$5101 N$5103 N$5212 N$5214 "Waveguide Crossing" sch_x=-118 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1373 N$5105 N$5107 N$5216 N$5218 "Waveguide Crossing" sch_x=-118 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1374 N$5109 N$5111 N$5220 N$5222 "Waveguide Crossing" sch_x=-118 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1375 N$5113 N$5115 N$5224 N$5226 "Waveguide Crossing" sch_x=-118 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1376 N$5117 N$5119 N$5228 N$5230 "Waveguide Crossing" sch_x=-118 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1377 N$5121 N$5123 N$5232 N$5234 "Waveguide Crossing" sch_x=-118 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1378 N$5125 N$5127 N$5236 N$5238 "Waveguide Crossing" sch_x=-118 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1379 N$5129 N$5131 N$5240 N$5242 "Waveguide Crossing" sch_x=-118 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1380 N$5133 N$5135 N$5244 N$5246 "Waveguide Crossing" sch_x=-118 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1381 N$5137 N$5139 N$5248 N$5250 "Waveguide Crossing" sch_x=-118 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1382 N$5141 N$5143 N$5252 N$5254 "Waveguide Crossing" sch_x=-118 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1383 N$5145 N$5147 N$5256 N$5258 "Waveguide Crossing" sch_x=-118 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1384 N$5149 N$5151 N$5260 N$5262 "Waveguide Crossing" sch_x=-118 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1385 N$5153 N$5155 N$5264 N$5266 "Waveguide Crossing" sch_x=-118 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1386 N$5157 N$5159 N$5268 N$5270 "Waveguide Crossing" sch_x=-118 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1387 N$5161 N$5163 N$5272 N$5274 "Waveguide Crossing" sch_x=-118 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1388 N$5165 N$5167 N$5276 N$5278 "Waveguide Crossing" sch_x=-118 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1389 N$5169 N$5171 N$5280 N$5282 "Waveguide Crossing" sch_x=-118 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1390 N$5173 N$5175 N$5284 N$5286 "Waveguide Crossing" sch_x=-118 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1391 N$5177 N$5179 N$5288 N$5290 "Waveguide Crossing" sch_x=-118 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1392 N$5181 N$5183 N$5292 N$5294 "Waveguide Crossing" sch_x=-118 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1393 N$5185 N$5187 N$5296 N$5298 "Waveguide Crossing" sch_x=-118 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1394 N$5189 N$5191 N$5300 N$5302 "Waveguide Crossing" sch_x=-118 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1395 N$5193 N$5195 N$5304 N$5306 "Waveguide Crossing" sch_x=-118 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1396 N$5197 N$5199 N$5308 N$5310 "Waveguide Crossing" sch_x=-118 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1397 N$5201 N$5203 N$5312 N$5314 "Waveguide Crossing" sch_x=-118 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1398 N$5205 N$5207 N$5316 N$6837 "Waveguide Crossing" sch_x=-118 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1399 N$5209 N$5211 N$6729 N$5318 "Waveguide Crossing" sch_x=-116 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1400 N$5213 N$5215 N$5320 N$5322 "Waveguide Crossing" sch_x=-116 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1401 N$5217 N$5219 N$5324 N$5326 "Waveguide Crossing" sch_x=-116 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1402 N$5221 N$5223 N$5328 N$5330 "Waveguide Crossing" sch_x=-116 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1403 N$5225 N$5227 N$5332 N$5334 "Waveguide Crossing" sch_x=-116 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1404 N$5229 N$5231 N$5336 N$5338 "Waveguide Crossing" sch_x=-116 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1405 N$5233 N$5235 N$5340 N$5342 "Waveguide Crossing" sch_x=-116 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1406 N$5237 N$5239 N$5344 N$5346 "Waveguide Crossing" sch_x=-116 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1407 N$5241 N$5243 N$5348 N$5350 "Waveguide Crossing" sch_x=-116 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1408 N$5245 N$5247 N$5352 N$5354 "Waveguide Crossing" sch_x=-116 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1409 N$5249 N$5251 N$5356 N$5358 "Waveguide Crossing" sch_x=-116 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1410 N$5253 N$5255 N$5360 N$5362 "Waveguide Crossing" sch_x=-116 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1411 N$5257 N$5259 N$5364 N$5366 "Waveguide Crossing" sch_x=-116 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1412 N$5261 N$5263 N$5368 N$5370 "Waveguide Crossing" sch_x=-116 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1413 N$5265 N$5267 N$5372 N$5374 "Waveguide Crossing" sch_x=-116 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1414 N$5269 N$5271 N$5376 N$5378 "Waveguide Crossing" sch_x=-116 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1415 N$5273 N$5275 N$5380 N$5382 "Waveguide Crossing" sch_x=-116 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1416 N$5277 N$5279 N$5384 N$5386 "Waveguide Crossing" sch_x=-116 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1417 N$5281 N$5283 N$5388 N$5390 "Waveguide Crossing" sch_x=-116 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1418 N$5285 N$5287 N$5392 N$5394 "Waveguide Crossing" sch_x=-116 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1419 N$5289 N$5291 N$5396 N$5398 "Waveguide Crossing" sch_x=-116 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1420 N$5293 N$5295 N$5400 N$5402 "Waveguide Crossing" sch_x=-116 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1421 N$5297 N$5299 N$5404 N$5406 "Waveguide Crossing" sch_x=-116 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1422 N$5301 N$5303 N$5408 N$5410 "Waveguide Crossing" sch_x=-116 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1423 N$5305 N$5307 N$5412 N$5414 "Waveguide Crossing" sch_x=-116 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1424 N$5309 N$5311 N$5416 N$5418 "Waveguide Crossing" sch_x=-116 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1425 N$5313 N$5315 N$5420 N$6835 "Waveguide Crossing" sch_x=-116 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1426 N$5317 N$5319 N$6731 N$5422 "Waveguide Crossing" sch_x=-114 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1427 N$5321 N$5323 N$5424 N$5426 "Waveguide Crossing" sch_x=-114 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1428 N$5325 N$5327 N$5428 N$5430 "Waveguide Crossing" sch_x=-114 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1429 N$5329 N$5331 N$5432 N$5434 "Waveguide Crossing" sch_x=-114 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1430 N$5333 N$5335 N$5436 N$5438 "Waveguide Crossing" sch_x=-114 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1431 N$5337 N$5339 N$5440 N$5442 "Waveguide Crossing" sch_x=-114 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1432 N$5341 N$5343 N$5444 N$5446 "Waveguide Crossing" sch_x=-114 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1433 N$5345 N$5347 N$5448 N$5450 "Waveguide Crossing" sch_x=-114 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1434 N$5349 N$5351 N$5452 N$5454 "Waveguide Crossing" sch_x=-114 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1435 N$5353 N$5355 N$5456 N$5458 "Waveguide Crossing" sch_x=-114 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1436 N$5357 N$5359 N$5460 N$5462 "Waveguide Crossing" sch_x=-114 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1437 N$5361 N$5363 N$5464 N$5466 "Waveguide Crossing" sch_x=-114 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1438 N$5365 N$5367 N$5468 N$5470 "Waveguide Crossing" sch_x=-114 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1439 N$5369 N$5371 N$5472 N$5474 "Waveguide Crossing" sch_x=-114 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1440 N$5373 N$5375 N$5476 N$5478 "Waveguide Crossing" sch_x=-114 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1441 N$5377 N$5379 N$5480 N$5482 "Waveguide Crossing" sch_x=-114 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1442 N$5381 N$5383 N$5484 N$5486 "Waveguide Crossing" sch_x=-114 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1443 N$5385 N$5387 N$5488 N$5490 "Waveguide Crossing" sch_x=-114 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1444 N$5389 N$5391 N$5492 N$5494 "Waveguide Crossing" sch_x=-114 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1445 N$5393 N$5395 N$5496 N$5498 "Waveguide Crossing" sch_x=-114 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1446 N$5397 N$5399 N$5500 N$5502 "Waveguide Crossing" sch_x=-114 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1447 N$5401 N$5403 N$5504 N$5506 "Waveguide Crossing" sch_x=-114 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1448 N$5405 N$5407 N$5508 N$5510 "Waveguide Crossing" sch_x=-114 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1449 N$5409 N$5411 N$5512 N$5514 "Waveguide Crossing" sch_x=-114 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1450 N$5413 N$5415 N$5516 N$5518 "Waveguide Crossing" sch_x=-114 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1451 N$5417 N$5419 N$5520 N$6833 "Waveguide Crossing" sch_x=-114 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1452 N$5421 N$5423 N$6733 N$5522 "Waveguide Crossing" sch_x=-112 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1453 N$5425 N$5427 N$5524 N$5526 "Waveguide Crossing" sch_x=-112 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1454 N$5429 N$5431 N$5528 N$5530 "Waveguide Crossing" sch_x=-112 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1455 N$5433 N$5435 N$5532 N$5534 "Waveguide Crossing" sch_x=-112 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1456 N$5437 N$5439 N$5536 N$5538 "Waveguide Crossing" sch_x=-112 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1457 N$5441 N$5443 N$5540 N$5542 "Waveguide Crossing" sch_x=-112 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1458 N$5445 N$5447 N$5544 N$5546 "Waveguide Crossing" sch_x=-112 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1459 N$5449 N$5451 N$5548 N$5550 "Waveguide Crossing" sch_x=-112 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1460 N$5453 N$5455 N$5552 N$5554 "Waveguide Crossing" sch_x=-112 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1461 N$5457 N$5459 N$5556 N$5558 "Waveguide Crossing" sch_x=-112 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1462 N$5461 N$5463 N$5560 N$5562 "Waveguide Crossing" sch_x=-112 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1463 N$5465 N$5467 N$5564 N$5566 "Waveguide Crossing" sch_x=-112 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1464 N$5469 N$5471 N$5568 N$5570 "Waveguide Crossing" sch_x=-112 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1465 N$5473 N$5475 N$5572 N$5574 "Waveguide Crossing" sch_x=-112 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1466 N$5477 N$5479 N$5576 N$5578 "Waveguide Crossing" sch_x=-112 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1467 N$5481 N$5483 N$5580 N$5582 "Waveguide Crossing" sch_x=-112 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1468 N$5485 N$5487 N$5584 N$5586 "Waveguide Crossing" sch_x=-112 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1469 N$5489 N$5491 N$5588 N$5590 "Waveguide Crossing" sch_x=-112 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1470 N$5493 N$5495 N$5592 N$5594 "Waveguide Crossing" sch_x=-112 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1471 N$5497 N$5499 N$5596 N$5598 "Waveguide Crossing" sch_x=-112 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1472 N$5501 N$5503 N$5600 N$5602 "Waveguide Crossing" sch_x=-112 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1473 N$5505 N$5507 N$5604 N$5606 "Waveguide Crossing" sch_x=-112 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1474 N$5509 N$5511 N$5608 N$5610 "Waveguide Crossing" sch_x=-112 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1475 N$5513 N$5515 N$5612 N$5614 "Waveguide Crossing" sch_x=-112 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1476 N$5517 N$5519 N$5616 N$6831 "Waveguide Crossing" sch_x=-112 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1477 N$5521 N$5523 N$6735 N$5618 "Waveguide Crossing" sch_x=-110 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1478 N$5525 N$5527 N$5620 N$5622 "Waveguide Crossing" sch_x=-110 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1479 N$5529 N$5531 N$5624 N$5626 "Waveguide Crossing" sch_x=-110 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1480 N$5533 N$5535 N$5628 N$5630 "Waveguide Crossing" sch_x=-110 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1481 N$5537 N$5539 N$5632 N$5634 "Waveguide Crossing" sch_x=-110 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1482 N$5541 N$5543 N$5636 N$5638 "Waveguide Crossing" sch_x=-110 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1483 N$5545 N$5547 N$5640 N$5642 "Waveguide Crossing" sch_x=-110 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1484 N$5549 N$5551 N$5644 N$5646 "Waveguide Crossing" sch_x=-110 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1485 N$5553 N$5555 N$5648 N$5650 "Waveguide Crossing" sch_x=-110 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1486 N$5557 N$5559 N$5652 N$5654 "Waveguide Crossing" sch_x=-110 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1487 N$5561 N$5563 N$5656 N$5658 "Waveguide Crossing" sch_x=-110 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1488 N$5565 N$5567 N$5660 N$5662 "Waveguide Crossing" sch_x=-110 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1489 N$5569 N$5571 N$5664 N$5666 "Waveguide Crossing" sch_x=-110 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1490 N$5573 N$5575 N$5668 N$5670 "Waveguide Crossing" sch_x=-110 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1491 N$5577 N$5579 N$5672 N$5674 "Waveguide Crossing" sch_x=-110 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1492 N$5581 N$5583 N$5676 N$5678 "Waveguide Crossing" sch_x=-110 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1493 N$5585 N$5587 N$5680 N$5682 "Waveguide Crossing" sch_x=-110 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1494 N$5589 N$5591 N$5684 N$5686 "Waveguide Crossing" sch_x=-110 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1495 N$5593 N$5595 N$5688 N$5690 "Waveguide Crossing" sch_x=-110 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1496 N$5597 N$5599 N$5692 N$5694 "Waveguide Crossing" sch_x=-110 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1497 N$5601 N$5603 N$5696 N$5698 "Waveguide Crossing" sch_x=-110 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1498 N$5605 N$5607 N$5700 N$5702 "Waveguide Crossing" sch_x=-110 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1499 N$5609 N$5611 N$5704 N$5706 "Waveguide Crossing" sch_x=-110 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1500 N$5613 N$5615 N$5708 N$6829 "Waveguide Crossing" sch_x=-110 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1501 N$5617 N$5619 N$6737 N$5710 "Waveguide Crossing" sch_x=-108 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1502 N$5621 N$5623 N$5712 N$5714 "Waveguide Crossing" sch_x=-108 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1503 N$5625 N$5627 N$5716 N$5718 "Waveguide Crossing" sch_x=-108 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1504 N$5629 N$5631 N$5720 N$5722 "Waveguide Crossing" sch_x=-108 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1505 N$5633 N$5635 N$5724 N$5726 "Waveguide Crossing" sch_x=-108 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1506 N$5637 N$5639 N$5728 N$5730 "Waveguide Crossing" sch_x=-108 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1507 N$5641 N$5643 N$5732 N$5734 "Waveguide Crossing" sch_x=-108 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1508 N$5645 N$5647 N$5736 N$5738 "Waveguide Crossing" sch_x=-108 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1509 N$5649 N$5651 N$5740 N$5742 "Waveguide Crossing" sch_x=-108 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1510 N$5653 N$5655 N$5744 N$5746 "Waveguide Crossing" sch_x=-108 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1511 N$5657 N$5659 N$5748 N$5750 "Waveguide Crossing" sch_x=-108 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1512 N$5661 N$5663 N$5752 N$5754 "Waveguide Crossing" sch_x=-108 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1513 N$5665 N$5667 N$5756 N$5758 "Waveguide Crossing" sch_x=-108 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1514 N$5669 N$5671 N$5760 N$5762 "Waveguide Crossing" sch_x=-108 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1515 N$5673 N$5675 N$5764 N$5766 "Waveguide Crossing" sch_x=-108 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1516 N$5677 N$5679 N$5768 N$5770 "Waveguide Crossing" sch_x=-108 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1517 N$5681 N$5683 N$5772 N$5774 "Waveguide Crossing" sch_x=-108 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1518 N$5685 N$5687 N$5776 N$5778 "Waveguide Crossing" sch_x=-108 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1519 N$5689 N$5691 N$5780 N$5782 "Waveguide Crossing" sch_x=-108 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1520 N$5693 N$5695 N$5784 N$5786 "Waveguide Crossing" sch_x=-108 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1521 N$5697 N$5699 N$5788 N$5790 "Waveguide Crossing" sch_x=-108 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1522 N$5701 N$5703 N$5792 N$5794 "Waveguide Crossing" sch_x=-108 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1523 N$5705 N$5707 N$5796 N$6827 "Waveguide Crossing" sch_x=-108 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1524 N$5709 N$5711 N$6739 N$5798 "Waveguide Crossing" sch_x=-106 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1525 N$5713 N$5715 N$5800 N$5802 "Waveguide Crossing" sch_x=-106 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1526 N$5717 N$5719 N$5804 N$5806 "Waveguide Crossing" sch_x=-106 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1527 N$5721 N$5723 N$5808 N$5810 "Waveguide Crossing" sch_x=-106 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1528 N$5725 N$5727 N$5812 N$5814 "Waveguide Crossing" sch_x=-106 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1529 N$5729 N$5731 N$5816 N$5818 "Waveguide Crossing" sch_x=-106 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1530 N$5733 N$5735 N$5820 N$5822 "Waveguide Crossing" sch_x=-106 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1531 N$5737 N$5739 N$5824 N$5826 "Waveguide Crossing" sch_x=-106 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1532 N$5741 N$5743 N$5828 N$5830 "Waveguide Crossing" sch_x=-106 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1533 N$5745 N$5747 N$5832 N$5834 "Waveguide Crossing" sch_x=-106 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1534 N$5749 N$5751 N$5836 N$5838 "Waveguide Crossing" sch_x=-106 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1535 N$5753 N$5755 N$5840 N$5842 "Waveguide Crossing" sch_x=-106 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1536 N$5757 N$5759 N$5844 N$5846 "Waveguide Crossing" sch_x=-106 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1537 N$5761 N$5763 N$5848 N$5850 "Waveguide Crossing" sch_x=-106 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1538 N$5765 N$5767 N$5852 N$5854 "Waveguide Crossing" sch_x=-106 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1539 N$5769 N$5771 N$5856 N$5858 "Waveguide Crossing" sch_x=-106 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1540 N$5773 N$5775 N$5860 N$5862 "Waveguide Crossing" sch_x=-106 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1541 N$5777 N$5779 N$5864 N$5866 "Waveguide Crossing" sch_x=-106 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1542 N$5781 N$5783 N$5868 N$5870 "Waveguide Crossing" sch_x=-106 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1543 N$5785 N$5787 N$5872 N$5874 "Waveguide Crossing" sch_x=-106 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1544 N$5789 N$5791 N$5876 N$5878 "Waveguide Crossing" sch_x=-106 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1545 N$5793 N$5795 N$5880 N$6825 "Waveguide Crossing" sch_x=-106 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1546 N$5797 N$5799 N$6741 N$5882 "Waveguide Crossing" sch_x=-104 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1547 N$5801 N$5803 N$5884 N$5886 "Waveguide Crossing" sch_x=-104 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1548 N$5805 N$5807 N$5888 N$5890 "Waveguide Crossing" sch_x=-104 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1549 N$5809 N$5811 N$5892 N$5894 "Waveguide Crossing" sch_x=-104 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1550 N$5813 N$5815 N$5896 N$5898 "Waveguide Crossing" sch_x=-104 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1551 N$5817 N$5819 N$5900 N$5902 "Waveguide Crossing" sch_x=-104 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1552 N$5821 N$5823 N$5904 N$5906 "Waveguide Crossing" sch_x=-104 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1553 N$5825 N$5827 N$5908 N$5910 "Waveguide Crossing" sch_x=-104 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1554 N$5829 N$5831 N$5912 N$5914 "Waveguide Crossing" sch_x=-104 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1555 N$5833 N$5835 N$5916 N$5918 "Waveguide Crossing" sch_x=-104 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1556 N$5837 N$5839 N$5920 N$5922 "Waveguide Crossing" sch_x=-104 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1557 N$5841 N$5843 N$5924 N$5926 "Waveguide Crossing" sch_x=-104 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1558 N$5845 N$5847 N$5928 N$5930 "Waveguide Crossing" sch_x=-104 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1559 N$5849 N$5851 N$5932 N$5934 "Waveguide Crossing" sch_x=-104 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1560 N$5853 N$5855 N$5936 N$5938 "Waveguide Crossing" sch_x=-104 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1561 N$5857 N$5859 N$5940 N$5942 "Waveguide Crossing" sch_x=-104 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1562 N$5861 N$5863 N$5944 N$5946 "Waveguide Crossing" sch_x=-104 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1563 N$5865 N$5867 N$5948 N$5950 "Waveguide Crossing" sch_x=-104 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1564 N$5869 N$5871 N$5952 N$5954 "Waveguide Crossing" sch_x=-104 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1565 N$5873 N$5875 N$5956 N$5958 "Waveguide Crossing" sch_x=-104 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1566 N$5877 N$5879 N$5960 N$6823 "Waveguide Crossing" sch_x=-104 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1567 N$5881 N$5883 N$6743 N$5962 "Waveguide Crossing" sch_x=-102 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1568 N$5885 N$5887 N$5964 N$5966 "Waveguide Crossing" sch_x=-102 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1569 N$5889 N$5891 N$5968 N$5970 "Waveguide Crossing" sch_x=-102 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1570 N$5893 N$5895 N$5972 N$5974 "Waveguide Crossing" sch_x=-102 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1571 N$5897 N$5899 N$5976 N$5978 "Waveguide Crossing" sch_x=-102 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1572 N$5901 N$5903 N$5980 N$5982 "Waveguide Crossing" sch_x=-102 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1573 N$5905 N$5907 N$5984 N$5986 "Waveguide Crossing" sch_x=-102 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1574 N$5909 N$5911 N$5988 N$5990 "Waveguide Crossing" sch_x=-102 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1575 N$5913 N$5915 N$5992 N$5994 "Waveguide Crossing" sch_x=-102 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1576 N$5917 N$5919 N$5996 N$5998 "Waveguide Crossing" sch_x=-102 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1577 N$5921 N$5923 N$6000 N$6002 "Waveguide Crossing" sch_x=-102 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1578 N$5925 N$5927 N$6004 N$6006 "Waveguide Crossing" sch_x=-102 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1579 N$5929 N$5931 N$6008 N$6010 "Waveguide Crossing" sch_x=-102 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1580 N$5933 N$5935 N$6012 N$6014 "Waveguide Crossing" sch_x=-102 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1581 N$5937 N$5939 N$6016 N$6018 "Waveguide Crossing" sch_x=-102 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1582 N$5941 N$5943 N$6020 N$6022 "Waveguide Crossing" sch_x=-102 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1583 N$5945 N$5947 N$6024 N$6026 "Waveguide Crossing" sch_x=-102 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1584 N$5949 N$5951 N$6028 N$6030 "Waveguide Crossing" sch_x=-102 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1585 N$5953 N$5955 N$6032 N$6034 "Waveguide Crossing" sch_x=-102 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1586 N$5957 N$5959 N$6036 N$6821 "Waveguide Crossing" sch_x=-102 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1587 N$5961 N$5963 N$6745 N$6038 "Waveguide Crossing" sch_x=-100 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1588 N$5965 N$5967 N$6040 N$6042 "Waveguide Crossing" sch_x=-100 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1589 N$5969 N$5971 N$6044 N$6046 "Waveguide Crossing" sch_x=-100 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1590 N$5973 N$5975 N$6048 N$6050 "Waveguide Crossing" sch_x=-100 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1591 N$5977 N$5979 N$6052 N$6054 "Waveguide Crossing" sch_x=-100 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1592 N$5981 N$5983 N$6056 N$6058 "Waveguide Crossing" sch_x=-100 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1593 N$5985 N$5987 N$6060 N$6062 "Waveguide Crossing" sch_x=-100 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1594 N$5989 N$5991 N$6064 N$6066 "Waveguide Crossing" sch_x=-100 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1595 N$5993 N$5995 N$6068 N$6070 "Waveguide Crossing" sch_x=-100 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1596 N$5997 N$5999 N$6072 N$6074 "Waveguide Crossing" sch_x=-100 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1597 N$6001 N$6003 N$6076 N$6078 "Waveguide Crossing" sch_x=-100 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1598 N$6005 N$6007 N$6080 N$6082 "Waveguide Crossing" sch_x=-100 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1599 N$6009 N$6011 N$6084 N$6086 "Waveguide Crossing" sch_x=-100 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1600 N$6013 N$6015 N$6088 N$6090 "Waveguide Crossing" sch_x=-100 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1601 N$6017 N$6019 N$6092 N$6094 "Waveguide Crossing" sch_x=-100 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1602 N$6021 N$6023 N$6096 N$6098 "Waveguide Crossing" sch_x=-100 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1603 N$6025 N$6027 N$6100 N$6102 "Waveguide Crossing" sch_x=-100 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1604 N$6029 N$6031 N$6104 N$6106 "Waveguide Crossing" sch_x=-100 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1605 N$6033 N$6035 N$6108 N$6819 "Waveguide Crossing" sch_x=-100 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1606 N$6037 N$6039 N$6747 N$6110 "Waveguide Crossing" sch_x=-98 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1607 N$6041 N$6043 N$6112 N$6114 "Waveguide Crossing" sch_x=-98 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1608 N$6045 N$6047 N$6116 N$6118 "Waveguide Crossing" sch_x=-98 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1609 N$6049 N$6051 N$6120 N$6122 "Waveguide Crossing" sch_x=-98 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1610 N$6053 N$6055 N$6124 N$6126 "Waveguide Crossing" sch_x=-98 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1611 N$6057 N$6059 N$6128 N$6130 "Waveguide Crossing" sch_x=-98 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1612 N$6061 N$6063 N$6132 N$6134 "Waveguide Crossing" sch_x=-98 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1613 N$6065 N$6067 N$6136 N$6138 "Waveguide Crossing" sch_x=-98 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1614 N$6069 N$6071 N$6140 N$6142 "Waveguide Crossing" sch_x=-98 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1615 N$6073 N$6075 N$6144 N$6146 "Waveguide Crossing" sch_x=-98 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1616 N$6077 N$6079 N$6148 N$6150 "Waveguide Crossing" sch_x=-98 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1617 N$6081 N$6083 N$6152 N$6154 "Waveguide Crossing" sch_x=-98 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1618 N$6085 N$6087 N$6156 N$6158 "Waveguide Crossing" sch_x=-98 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1619 N$6089 N$6091 N$6160 N$6162 "Waveguide Crossing" sch_x=-98 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1620 N$6093 N$6095 N$6164 N$6166 "Waveguide Crossing" sch_x=-98 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1621 N$6097 N$6099 N$6168 N$6170 "Waveguide Crossing" sch_x=-98 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1622 N$6101 N$6103 N$6172 N$6174 "Waveguide Crossing" sch_x=-98 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1623 N$6105 N$6107 N$6176 N$6817 "Waveguide Crossing" sch_x=-98 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1624 N$6109 N$6111 N$6749 N$6178 "Waveguide Crossing" sch_x=-96 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1625 N$6113 N$6115 N$6180 N$6182 "Waveguide Crossing" sch_x=-96 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1626 N$6117 N$6119 N$6184 N$6186 "Waveguide Crossing" sch_x=-96 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1627 N$6121 N$6123 N$6188 N$6190 "Waveguide Crossing" sch_x=-96 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1628 N$6125 N$6127 N$6192 N$6194 "Waveguide Crossing" sch_x=-96 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1629 N$6129 N$6131 N$6196 N$6198 "Waveguide Crossing" sch_x=-96 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1630 N$6133 N$6135 N$6200 N$6202 "Waveguide Crossing" sch_x=-96 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1631 N$6137 N$6139 N$6204 N$6206 "Waveguide Crossing" sch_x=-96 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1632 N$6141 N$6143 N$6208 N$6210 "Waveguide Crossing" sch_x=-96 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1633 N$6145 N$6147 N$6212 N$6214 "Waveguide Crossing" sch_x=-96 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1634 N$6149 N$6151 N$6216 N$6218 "Waveguide Crossing" sch_x=-96 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1635 N$6153 N$6155 N$6220 N$6222 "Waveguide Crossing" sch_x=-96 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1636 N$6157 N$6159 N$6224 N$6226 "Waveguide Crossing" sch_x=-96 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1637 N$6161 N$6163 N$6228 N$6230 "Waveguide Crossing" sch_x=-96 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1638 N$6165 N$6167 N$6232 N$6234 "Waveguide Crossing" sch_x=-96 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1639 N$6169 N$6171 N$6236 N$6238 "Waveguide Crossing" sch_x=-96 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1640 N$6173 N$6175 N$6240 N$6815 "Waveguide Crossing" sch_x=-96 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1641 N$6177 N$6179 N$6751 N$6242 "Waveguide Crossing" sch_x=-94 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1642 N$6181 N$6183 N$6244 N$6246 "Waveguide Crossing" sch_x=-94 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1643 N$6185 N$6187 N$6248 N$6250 "Waveguide Crossing" sch_x=-94 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1644 N$6189 N$6191 N$6252 N$6254 "Waveguide Crossing" sch_x=-94 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1645 N$6193 N$6195 N$6256 N$6258 "Waveguide Crossing" sch_x=-94 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1646 N$6197 N$6199 N$6260 N$6262 "Waveguide Crossing" sch_x=-94 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1647 N$6201 N$6203 N$6264 N$6266 "Waveguide Crossing" sch_x=-94 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1648 N$6205 N$6207 N$6268 N$6270 "Waveguide Crossing" sch_x=-94 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1649 N$6209 N$6211 N$6272 N$6274 "Waveguide Crossing" sch_x=-94 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1650 N$6213 N$6215 N$6276 N$6278 "Waveguide Crossing" sch_x=-94 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1651 N$6217 N$6219 N$6280 N$6282 "Waveguide Crossing" sch_x=-94 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1652 N$6221 N$6223 N$6284 N$6286 "Waveguide Crossing" sch_x=-94 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1653 N$6225 N$6227 N$6288 N$6290 "Waveguide Crossing" sch_x=-94 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1654 N$6229 N$6231 N$6292 N$6294 "Waveguide Crossing" sch_x=-94 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1655 N$6233 N$6235 N$6296 N$6298 "Waveguide Crossing" sch_x=-94 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1656 N$6237 N$6239 N$6300 N$6813 "Waveguide Crossing" sch_x=-94 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1657 N$6241 N$6243 N$6753 N$6302 "Waveguide Crossing" sch_x=-92 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1658 N$6245 N$6247 N$6304 N$6306 "Waveguide Crossing" sch_x=-92 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1659 N$6249 N$6251 N$6308 N$6310 "Waveguide Crossing" sch_x=-92 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1660 N$6253 N$6255 N$6312 N$6314 "Waveguide Crossing" sch_x=-92 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1661 N$6257 N$6259 N$6316 N$6318 "Waveguide Crossing" sch_x=-92 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1662 N$6261 N$6263 N$6320 N$6322 "Waveguide Crossing" sch_x=-92 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1663 N$6265 N$6267 N$6324 N$6326 "Waveguide Crossing" sch_x=-92 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1664 N$6269 N$6271 N$6328 N$6330 "Waveguide Crossing" sch_x=-92 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1665 N$6273 N$6275 N$6332 N$6334 "Waveguide Crossing" sch_x=-92 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1666 N$6277 N$6279 N$6336 N$6338 "Waveguide Crossing" sch_x=-92 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1667 N$6281 N$6283 N$6340 N$6342 "Waveguide Crossing" sch_x=-92 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1668 N$6285 N$6287 N$6344 N$6346 "Waveguide Crossing" sch_x=-92 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1669 N$6289 N$6291 N$6348 N$6350 "Waveguide Crossing" sch_x=-92 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1670 N$6293 N$6295 N$6352 N$6354 "Waveguide Crossing" sch_x=-92 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1671 N$6297 N$6299 N$6356 N$6811 "Waveguide Crossing" sch_x=-92 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1672 N$6301 N$6303 N$6755 N$6358 "Waveguide Crossing" sch_x=-90 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1673 N$6305 N$6307 N$6360 N$6362 "Waveguide Crossing" sch_x=-90 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1674 N$6309 N$6311 N$6364 N$6366 "Waveguide Crossing" sch_x=-90 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1675 N$6313 N$6315 N$6368 N$6370 "Waveguide Crossing" sch_x=-90 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1676 N$6317 N$6319 N$6372 N$6374 "Waveguide Crossing" sch_x=-90 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1677 N$6321 N$6323 N$6376 N$6378 "Waveguide Crossing" sch_x=-90 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1678 N$6325 N$6327 N$6380 N$6382 "Waveguide Crossing" sch_x=-90 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1679 N$6329 N$6331 N$6384 N$6386 "Waveguide Crossing" sch_x=-90 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1680 N$6333 N$6335 N$6388 N$6390 "Waveguide Crossing" sch_x=-90 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1681 N$6337 N$6339 N$6392 N$6394 "Waveguide Crossing" sch_x=-90 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1682 N$6341 N$6343 N$6396 N$6398 "Waveguide Crossing" sch_x=-90 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1683 N$6345 N$6347 N$6400 N$6402 "Waveguide Crossing" sch_x=-90 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1684 N$6349 N$6351 N$6404 N$6406 "Waveguide Crossing" sch_x=-90 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1685 N$6353 N$6355 N$6408 N$6809 "Waveguide Crossing" sch_x=-90 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1686 N$6357 N$6359 N$6757 N$6410 "Waveguide Crossing" sch_x=-88 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1687 N$6361 N$6363 N$6412 N$6414 "Waveguide Crossing" sch_x=-88 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1688 N$6365 N$6367 N$6416 N$6418 "Waveguide Crossing" sch_x=-88 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1689 N$6369 N$6371 N$6420 N$6422 "Waveguide Crossing" sch_x=-88 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1690 N$6373 N$6375 N$6424 N$6426 "Waveguide Crossing" sch_x=-88 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1691 N$6377 N$6379 N$6428 N$6430 "Waveguide Crossing" sch_x=-88 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1692 N$6381 N$6383 N$6432 N$6434 "Waveguide Crossing" sch_x=-88 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1693 N$6385 N$6387 N$6436 N$6438 "Waveguide Crossing" sch_x=-88 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1694 N$6389 N$6391 N$6440 N$6442 "Waveguide Crossing" sch_x=-88 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1695 N$6393 N$6395 N$6444 N$6446 "Waveguide Crossing" sch_x=-88 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1696 N$6397 N$6399 N$6448 N$6450 "Waveguide Crossing" sch_x=-88 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1697 N$6401 N$6403 N$6452 N$6454 "Waveguide Crossing" sch_x=-88 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1698 N$6405 N$6407 N$6456 N$6807 "Waveguide Crossing" sch_x=-88 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1699 N$6409 N$6411 N$6759 N$6458 "Waveguide Crossing" sch_x=-86 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1700 N$6413 N$6415 N$6460 N$6462 "Waveguide Crossing" sch_x=-86 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1701 N$6417 N$6419 N$6464 N$6466 "Waveguide Crossing" sch_x=-86 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1702 N$6421 N$6423 N$6468 N$6470 "Waveguide Crossing" sch_x=-86 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1703 N$6425 N$6427 N$6472 N$6474 "Waveguide Crossing" sch_x=-86 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1704 N$6429 N$6431 N$6476 N$6478 "Waveguide Crossing" sch_x=-86 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1705 N$6433 N$6435 N$6480 N$6482 "Waveguide Crossing" sch_x=-86 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1706 N$6437 N$6439 N$6484 N$6486 "Waveguide Crossing" sch_x=-86 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1707 N$6441 N$6443 N$6488 N$6490 "Waveguide Crossing" sch_x=-86 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1708 N$6445 N$6447 N$6492 N$6494 "Waveguide Crossing" sch_x=-86 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1709 N$6449 N$6451 N$6496 N$6498 "Waveguide Crossing" sch_x=-86 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1710 N$6453 N$6455 N$6500 N$6805 "Waveguide Crossing" sch_x=-86 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1711 N$6457 N$6459 N$6761 N$6502 "Waveguide Crossing" sch_x=-84 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1712 N$6461 N$6463 N$6504 N$6506 "Waveguide Crossing" sch_x=-84 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1713 N$6465 N$6467 N$6508 N$6510 "Waveguide Crossing" sch_x=-84 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1714 N$6469 N$6471 N$6512 N$6514 "Waveguide Crossing" sch_x=-84 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1715 N$6473 N$6475 N$6516 N$6518 "Waveguide Crossing" sch_x=-84 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1716 N$6477 N$6479 N$6520 N$6522 "Waveguide Crossing" sch_x=-84 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1717 N$6481 N$6483 N$6524 N$6526 "Waveguide Crossing" sch_x=-84 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1718 N$6485 N$6487 N$6528 N$6530 "Waveguide Crossing" sch_x=-84 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1719 N$6489 N$6491 N$6532 N$6534 "Waveguide Crossing" sch_x=-84 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1720 N$6493 N$6495 N$6536 N$6538 "Waveguide Crossing" sch_x=-84 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1721 N$6497 N$6499 N$6540 N$6803 "Waveguide Crossing" sch_x=-84 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1722 N$6501 N$6503 N$6763 N$6542 "Waveguide Crossing" sch_x=-82 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1723 N$6505 N$6507 N$6544 N$6546 "Waveguide Crossing" sch_x=-82 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1724 N$6509 N$6511 N$6548 N$6550 "Waveguide Crossing" sch_x=-82 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1725 N$6513 N$6515 N$6552 N$6554 "Waveguide Crossing" sch_x=-82 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1726 N$6517 N$6519 N$6556 N$6558 "Waveguide Crossing" sch_x=-82 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1727 N$6521 N$6523 N$6560 N$6562 "Waveguide Crossing" sch_x=-82 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1728 N$6525 N$6527 N$6564 N$6566 "Waveguide Crossing" sch_x=-82 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1729 N$6529 N$6531 N$6568 N$6570 "Waveguide Crossing" sch_x=-82 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1730 N$6533 N$6535 N$6572 N$6574 "Waveguide Crossing" sch_x=-82 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1731 N$6537 N$6539 N$6576 N$6801 "Waveguide Crossing" sch_x=-82 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1732 N$6541 N$6543 N$6765 N$6578 "Waveguide Crossing" sch_x=-80 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1733 N$6545 N$6547 N$6580 N$6582 "Waveguide Crossing" sch_x=-80 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1734 N$6549 N$6551 N$6584 N$6586 "Waveguide Crossing" sch_x=-80 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1735 N$6553 N$6555 N$6588 N$6590 "Waveguide Crossing" sch_x=-80 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1736 N$6557 N$6559 N$6592 N$6594 "Waveguide Crossing" sch_x=-80 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1737 N$6561 N$6563 N$6596 N$6598 "Waveguide Crossing" sch_x=-80 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1738 N$6565 N$6567 N$6600 N$6602 "Waveguide Crossing" sch_x=-80 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1739 N$6569 N$6571 N$6604 N$6606 "Waveguide Crossing" sch_x=-80 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1740 N$6573 N$6575 N$6608 N$6799 "Waveguide Crossing" sch_x=-80 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1741 N$6577 N$6579 N$6767 N$6610 "Waveguide Crossing" sch_x=-78 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1742 N$6581 N$6583 N$6612 N$6614 "Waveguide Crossing" sch_x=-78 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1743 N$6585 N$6587 N$6616 N$6618 "Waveguide Crossing" sch_x=-78 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1744 N$6589 N$6591 N$6620 N$6622 "Waveguide Crossing" sch_x=-78 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1745 N$6593 N$6595 N$6624 N$6626 "Waveguide Crossing" sch_x=-78 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1746 N$6597 N$6599 N$6628 N$6630 "Waveguide Crossing" sch_x=-78 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1747 N$6601 N$6603 N$6632 N$6634 "Waveguide Crossing" sch_x=-78 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1748 N$6605 N$6607 N$6636 N$6797 "Waveguide Crossing" sch_x=-78 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1749 N$6609 N$6611 N$6769 N$6638 "Waveguide Crossing" sch_x=-76 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1750 N$6613 N$6615 N$6640 N$6642 "Waveguide Crossing" sch_x=-76 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1751 N$6617 N$6619 N$6644 N$6646 "Waveguide Crossing" sch_x=-76 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1752 N$6621 N$6623 N$6648 N$6650 "Waveguide Crossing" sch_x=-76 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1753 N$6625 N$6627 N$6652 N$6654 "Waveguide Crossing" sch_x=-76 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1754 N$6629 N$6631 N$6656 N$6658 "Waveguide Crossing" sch_x=-76 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1755 N$6633 N$6635 N$6660 N$6795 "Waveguide Crossing" sch_x=-76 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1756 N$6637 N$6639 N$6771 N$6662 "Waveguide Crossing" sch_x=-74 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1757 N$6641 N$6643 N$6664 N$6666 "Waveguide Crossing" sch_x=-74 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1758 N$6645 N$6647 N$6668 N$6670 "Waveguide Crossing" sch_x=-74 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1759 N$6649 N$6651 N$6672 N$6674 "Waveguide Crossing" sch_x=-74 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1760 N$6653 N$6655 N$6676 N$6678 "Waveguide Crossing" sch_x=-74 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1761 N$6657 N$6659 N$6680 N$6793 "Waveguide Crossing" sch_x=-74 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1762 N$6661 N$6663 N$6773 N$6682 "Waveguide Crossing" sch_x=-72 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1763 N$6665 N$6667 N$6684 N$6686 "Waveguide Crossing" sch_x=-72 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1764 N$6669 N$6671 N$6688 N$6690 "Waveguide Crossing" sch_x=-72 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1765 N$6673 N$6675 N$6692 N$6694 "Waveguide Crossing" sch_x=-72 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1766 N$6677 N$6679 N$6696 N$6791 "Waveguide Crossing" sch_x=-72 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1767 N$6681 N$6683 N$6775 N$6698 "Waveguide Crossing" sch_x=-70 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1768 N$6685 N$6687 N$6700 N$6702 "Waveguide Crossing" sch_x=-70 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1769 N$6689 N$6691 N$6704 N$6706 "Waveguide Crossing" sch_x=-70 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1770 N$6693 N$6695 N$6708 N$6789 "Waveguide Crossing" sch_x=-70 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1771 N$6697 N$6699 N$6777 N$6710 "Waveguide Crossing" sch_x=-68 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1772 N$6701 N$6703 N$6712 N$6714 "Waveguide Crossing" sch_x=-68 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1773 N$6705 N$6707 N$6716 N$6787 "Waveguide Crossing" sch_x=-68 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1774 N$6709 N$6711 N$6779 N$6718 "Waveguide Crossing" sch_x=-66 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1775 N$6713 N$6715 N$6720 N$6785 "Waveguide Crossing" sch_x=-66 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1776 N$6717 N$6719 N$6781 N$6783 "Waveguide Crossing" sch_x=-64 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S977 N$6784 N$6786 N$4189 N$3650 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S978 N$6788 N$6790 N$3652 N$3654 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S979 N$6792 N$6794 N$3656 N$3658 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S980 N$6796 N$6798 N$3660 N$3662 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S981 N$6800 N$6802 N$3664 N$3666 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S982 N$6804 N$6806 N$3668 N$3670 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S983 N$6808 N$6810 N$3672 N$3674 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S984 N$6812 N$6814 N$3676 N$3678 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S985 N$6816 N$6818 N$3680 N$3682 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S986 N$6820 N$6822 N$3684 N$3686 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S987 N$6824 N$6826 N$3688 N$3690 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S988 N$6828 N$6830 N$3692 N$3694 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S989 N$6832 N$6834 N$3696 N$3698 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S990 N$6836 N$6838 N$3700 N$3702 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S991 N$6840 N$6842 N$3704 N$3706 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S992 N$6844 N$6848 N$3708 N$4191 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C993 N$3649 N$3651 N$4129 N$3710 "Waveguide Crossing" sch_x=-60 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C994 N$3653 N$3655 N$3712 N$3714 "Waveguide Crossing" sch_x=-60 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C995 N$3657 N$3659 N$3716 N$3718 "Waveguide Crossing" sch_x=-60 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C996 N$3661 N$3663 N$3720 N$3722 "Waveguide Crossing" sch_x=-60 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C997 N$3665 N$3667 N$3724 N$3726 "Waveguide Crossing" sch_x=-60 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C998 N$3669 N$3671 N$3728 N$3730 "Waveguide Crossing" sch_x=-60 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C999 N$3673 N$3675 N$3732 N$3734 "Waveguide Crossing" sch_x=-60 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1000 N$3677 N$3679 N$3736 N$3738 "Waveguide Crossing" sch_x=-60 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1001 N$3681 N$3683 N$3740 N$3742 "Waveguide Crossing" sch_x=-60 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1002 N$3685 N$3687 N$3744 N$3746 "Waveguide Crossing" sch_x=-60 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1003 N$3689 N$3691 N$3748 N$3750 "Waveguide Crossing" sch_x=-60 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1004 N$3693 N$3695 N$3752 N$3754 "Waveguide Crossing" sch_x=-60 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1005 N$3697 N$3699 N$3756 N$3758 "Waveguide Crossing" sch_x=-60 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1006 N$3701 N$3703 N$3760 N$3762 "Waveguide Crossing" sch_x=-60 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1007 N$3705 N$3707 N$3764 N$4187 "Waveguide Crossing" sch_x=-60 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1008 N$3709 N$3711 N$4131 N$3766 "Waveguide Crossing" sch_x=-58 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1009 N$3713 N$3715 N$3768 N$3770 "Waveguide Crossing" sch_x=-58 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1010 N$3717 N$3719 N$3772 N$3774 "Waveguide Crossing" sch_x=-58 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1011 N$3721 N$3723 N$3776 N$3778 "Waveguide Crossing" sch_x=-58 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1012 N$3725 N$3727 N$3780 N$3782 "Waveguide Crossing" sch_x=-58 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1013 N$3729 N$3731 N$3784 N$3786 "Waveguide Crossing" sch_x=-58 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1014 N$3733 N$3735 N$3788 N$3790 "Waveguide Crossing" sch_x=-58 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1015 N$3737 N$3739 N$3792 N$3794 "Waveguide Crossing" sch_x=-58 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1016 N$3741 N$3743 N$3796 N$3798 "Waveguide Crossing" sch_x=-58 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1017 N$3745 N$3747 N$3800 N$3802 "Waveguide Crossing" sch_x=-58 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1018 N$3749 N$3751 N$3804 N$3806 "Waveguide Crossing" sch_x=-58 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1019 N$3753 N$3755 N$3808 N$3810 "Waveguide Crossing" sch_x=-58 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1020 N$3757 N$3759 N$3812 N$3814 "Waveguide Crossing" sch_x=-58 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1021 N$3761 N$3763 N$3816 N$4185 "Waveguide Crossing" sch_x=-58 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1022 N$3765 N$3767 N$4133 N$3818 "Waveguide Crossing" sch_x=-56 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1023 N$3769 N$3771 N$3820 N$3822 "Waveguide Crossing" sch_x=-56 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1024 N$3773 N$3775 N$3824 N$3826 "Waveguide Crossing" sch_x=-56 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1025 N$3777 N$3779 N$3828 N$3830 "Waveguide Crossing" sch_x=-56 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1026 N$3781 N$3783 N$3832 N$3834 "Waveguide Crossing" sch_x=-56 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1027 N$3785 N$3787 N$3836 N$3838 "Waveguide Crossing" sch_x=-56 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1028 N$3789 N$3791 N$3840 N$3842 "Waveguide Crossing" sch_x=-56 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1029 N$3793 N$3795 N$3844 N$3846 "Waveguide Crossing" sch_x=-56 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1030 N$3797 N$3799 N$3848 N$3850 "Waveguide Crossing" sch_x=-56 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1031 N$3801 N$3803 N$3852 N$3854 "Waveguide Crossing" sch_x=-56 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1032 N$3805 N$3807 N$3856 N$3858 "Waveguide Crossing" sch_x=-56 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1033 N$3809 N$3811 N$3860 N$3862 "Waveguide Crossing" sch_x=-56 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1034 N$3813 N$3815 N$3864 N$4183 "Waveguide Crossing" sch_x=-56 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1035 N$3817 N$3819 N$4135 N$3866 "Waveguide Crossing" sch_x=-54 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1036 N$3821 N$3823 N$3868 N$3870 "Waveguide Crossing" sch_x=-54 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1037 N$3825 N$3827 N$3872 N$3874 "Waveguide Crossing" sch_x=-54 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1038 N$3829 N$3831 N$3876 N$3878 "Waveguide Crossing" sch_x=-54 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1039 N$3833 N$3835 N$3880 N$3882 "Waveguide Crossing" sch_x=-54 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1040 N$3837 N$3839 N$3884 N$3886 "Waveguide Crossing" sch_x=-54 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1041 N$3841 N$3843 N$3888 N$3890 "Waveguide Crossing" sch_x=-54 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1042 N$3845 N$3847 N$3892 N$3894 "Waveguide Crossing" sch_x=-54 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1043 N$3849 N$3851 N$3896 N$3898 "Waveguide Crossing" sch_x=-54 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1044 N$3853 N$3855 N$3900 N$3902 "Waveguide Crossing" sch_x=-54 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1045 N$3857 N$3859 N$3904 N$3906 "Waveguide Crossing" sch_x=-54 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1046 N$3861 N$3863 N$3908 N$4181 "Waveguide Crossing" sch_x=-54 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1047 N$3865 N$3867 N$4137 N$3910 "Waveguide Crossing" sch_x=-52 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1048 N$3869 N$3871 N$3912 N$3914 "Waveguide Crossing" sch_x=-52 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1049 N$3873 N$3875 N$3916 N$3918 "Waveguide Crossing" sch_x=-52 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1050 N$3877 N$3879 N$3920 N$3922 "Waveguide Crossing" sch_x=-52 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1051 N$3881 N$3883 N$3924 N$3926 "Waveguide Crossing" sch_x=-52 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1052 N$3885 N$3887 N$3928 N$3930 "Waveguide Crossing" sch_x=-52 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1053 N$3889 N$3891 N$3932 N$3934 "Waveguide Crossing" sch_x=-52 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1054 N$3893 N$3895 N$3936 N$3938 "Waveguide Crossing" sch_x=-52 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1055 N$3897 N$3899 N$3940 N$3942 "Waveguide Crossing" sch_x=-52 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1056 N$3901 N$3903 N$3944 N$3946 "Waveguide Crossing" sch_x=-52 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1057 N$3905 N$3907 N$3948 N$4179 "Waveguide Crossing" sch_x=-52 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1058 N$3909 N$3911 N$4139 N$3950 "Waveguide Crossing" sch_x=-50 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1059 N$3913 N$3915 N$3952 N$3954 "Waveguide Crossing" sch_x=-50 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1060 N$3917 N$3919 N$3956 N$3958 "Waveguide Crossing" sch_x=-50 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1061 N$3921 N$3923 N$3960 N$3962 "Waveguide Crossing" sch_x=-50 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1062 N$3925 N$3927 N$3964 N$3966 "Waveguide Crossing" sch_x=-50 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1063 N$3929 N$3931 N$3968 N$3970 "Waveguide Crossing" sch_x=-50 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1064 N$3933 N$3935 N$3972 N$3974 "Waveguide Crossing" sch_x=-50 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1065 N$3937 N$3939 N$3976 N$3978 "Waveguide Crossing" sch_x=-50 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1066 N$3941 N$3943 N$3980 N$3982 "Waveguide Crossing" sch_x=-50 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1067 N$3945 N$3947 N$3984 N$4177 "Waveguide Crossing" sch_x=-50 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1068 N$3949 N$3951 N$4141 N$3986 "Waveguide Crossing" sch_x=-48 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1069 N$3953 N$3955 N$3988 N$3990 "Waveguide Crossing" sch_x=-48 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1070 N$3957 N$3959 N$3992 N$3994 "Waveguide Crossing" sch_x=-48 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1071 N$3961 N$3963 N$3996 N$3998 "Waveguide Crossing" sch_x=-48 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1072 N$3965 N$3967 N$4000 N$4002 "Waveguide Crossing" sch_x=-48 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1073 N$3969 N$3971 N$4004 N$4006 "Waveguide Crossing" sch_x=-48 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1074 N$3973 N$3975 N$4008 N$4010 "Waveguide Crossing" sch_x=-48 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1075 N$3977 N$3979 N$4012 N$4014 "Waveguide Crossing" sch_x=-48 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1076 N$3981 N$3983 N$4016 N$4175 "Waveguide Crossing" sch_x=-48 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1077 N$3985 N$3987 N$4143 N$4018 "Waveguide Crossing" sch_x=-46 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1078 N$3989 N$3991 N$4020 N$4022 "Waveguide Crossing" sch_x=-46 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1079 N$3993 N$3995 N$4024 N$4026 "Waveguide Crossing" sch_x=-46 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1080 N$3997 N$3999 N$4028 N$4030 "Waveguide Crossing" sch_x=-46 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1081 N$4001 N$4003 N$4032 N$4034 "Waveguide Crossing" sch_x=-46 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1082 N$4005 N$4007 N$4036 N$4038 "Waveguide Crossing" sch_x=-46 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1083 N$4009 N$4011 N$4040 N$4042 "Waveguide Crossing" sch_x=-46 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1084 N$4013 N$4015 N$4044 N$4173 "Waveguide Crossing" sch_x=-46 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1085 N$4017 N$4019 N$4145 N$4046 "Waveguide Crossing" sch_x=-44 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1086 N$4021 N$4023 N$4048 N$4050 "Waveguide Crossing" sch_x=-44 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1087 N$4025 N$4027 N$4052 N$4054 "Waveguide Crossing" sch_x=-44 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1088 N$4029 N$4031 N$4056 N$4058 "Waveguide Crossing" sch_x=-44 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1089 N$4033 N$4035 N$4060 N$4062 "Waveguide Crossing" sch_x=-44 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1090 N$4037 N$4039 N$4064 N$4066 "Waveguide Crossing" sch_x=-44 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1091 N$4041 N$4043 N$4068 N$4171 "Waveguide Crossing" sch_x=-44 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1092 N$4045 N$4047 N$4147 N$4070 "Waveguide Crossing" sch_x=-42 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1093 N$4049 N$4051 N$4072 N$4074 "Waveguide Crossing" sch_x=-42 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1094 N$4053 N$4055 N$4076 N$4078 "Waveguide Crossing" sch_x=-42 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1095 N$4057 N$4059 N$4080 N$4082 "Waveguide Crossing" sch_x=-42 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1096 N$4061 N$4063 N$4084 N$4086 "Waveguide Crossing" sch_x=-42 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1097 N$4065 N$4067 N$4088 N$4169 "Waveguide Crossing" sch_x=-42 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1098 N$4069 N$4071 N$4149 N$4090 "Waveguide Crossing" sch_x=-40 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1099 N$4073 N$4075 N$4092 N$4094 "Waveguide Crossing" sch_x=-40 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1100 N$4077 N$4079 N$4096 N$4098 "Waveguide Crossing" sch_x=-40 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1101 N$4081 N$4083 N$4100 N$4102 "Waveguide Crossing" sch_x=-40 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1102 N$4085 N$4087 N$4104 N$4167 "Waveguide Crossing" sch_x=-40 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1103 N$4089 N$4091 N$4151 N$4106 "Waveguide Crossing" sch_x=-38 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1104 N$4093 N$4095 N$4108 N$4110 "Waveguide Crossing" sch_x=-38 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1105 N$4097 N$4099 N$4112 N$4114 "Waveguide Crossing" sch_x=-38 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1106 N$4101 N$4103 N$4116 N$4165 "Waveguide Crossing" sch_x=-38 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1107 N$4105 N$4107 N$4153 N$4118 "Waveguide Crossing" sch_x=-36 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1108 N$4109 N$4111 N$4120 N$4122 "Waveguide Crossing" sch_x=-36 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1109 N$4113 N$4115 N$4124 N$4163 "Waveguide Crossing" sch_x=-36 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1110 N$4117 N$4119 N$4155 N$4126 "Waveguide Crossing" sch_x=-34 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1111 N$4121 N$4123 N$4128 N$4161 "Waveguide Crossing" sch_x=-34 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1112 N$4125 N$4127 N$4157 N$4159 "Waveguide Crossing" sch_x=-32 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S905 N$4160 N$4162 N$3501 N$3362 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S906 N$4164 N$4166 N$3364 N$3366 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S907 N$4168 N$4170 N$3368 N$3370 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S908 N$4172 N$4174 N$3372 N$3374 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S909 N$4176 N$4178 N$3376 N$3378 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S910 N$4180 N$4182 N$3380 N$3382 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S911 N$4184 N$4186 N$3384 N$3386 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S912 N$4188 N$4192 N$3388 N$3503 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C913 N$3361 N$3363 N$3473 N$3390 "Waveguide Crossing" sch_x=-28 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C914 N$3365 N$3367 N$3392 N$3394 "Waveguide Crossing" sch_x=-28 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C915 N$3369 N$3371 N$3396 N$3398 "Waveguide Crossing" sch_x=-28 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C916 N$3373 N$3375 N$3400 N$3402 "Waveguide Crossing" sch_x=-28 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C917 N$3377 N$3379 N$3404 N$3406 "Waveguide Crossing" sch_x=-28 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C918 N$3381 N$3383 N$3408 N$3410 "Waveguide Crossing" sch_x=-28 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C919 N$3385 N$3387 N$3412 N$3499 "Waveguide Crossing" sch_x=-28 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C920 N$3389 N$3391 N$3475 N$3414 "Waveguide Crossing" sch_x=-26 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C921 N$3393 N$3395 N$3416 N$3418 "Waveguide Crossing" sch_x=-26 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C922 N$3397 N$3399 N$3420 N$3422 "Waveguide Crossing" sch_x=-26 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C923 N$3401 N$3403 N$3424 N$3426 "Waveguide Crossing" sch_x=-26 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C924 N$3405 N$3407 N$3428 N$3430 "Waveguide Crossing" sch_x=-26 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C925 N$3409 N$3411 N$3432 N$3497 "Waveguide Crossing" sch_x=-26 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C926 N$3413 N$3415 N$3477 N$3434 "Waveguide Crossing" sch_x=-24 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C927 N$3417 N$3419 N$3436 N$3438 "Waveguide Crossing" sch_x=-24 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C928 N$3421 N$3423 N$3440 N$3442 "Waveguide Crossing" sch_x=-24 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C929 N$3425 N$3427 N$3444 N$3446 "Waveguide Crossing" sch_x=-24 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C930 N$3429 N$3431 N$3448 N$3495 "Waveguide Crossing" sch_x=-24 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C931 N$3433 N$3435 N$3479 N$3450 "Waveguide Crossing" sch_x=-22 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C932 N$3437 N$3439 N$3452 N$3454 "Waveguide Crossing" sch_x=-22 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C933 N$3441 N$3443 N$3456 N$3458 "Waveguide Crossing" sch_x=-22 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C934 N$3445 N$3447 N$3460 N$3493 "Waveguide Crossing" sch_x=-22 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C935 N$3449 N$3451 N$3481 N$3462 "Waveguide Crossing" sch_x=-20 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C936 N$3453 N$3455 N$3464 N$3466 "Waveguide Crossing" sch_x=-20 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C937 N$3457 N$3459 N$3468 N$3491 "Waveguide Crossing" sch_x=-20 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C938 N$3461 N$3463 N$3483 N$3470 "Waveguide Crossing" sch_x=-18 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C939 N$3465 N$3467 N$3472 N$3489 "Waveguide Crossing" sch_x=-18 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C940 N$3469 N$3471 N$3485 N$3487 "Waveguide Crossing" sch_x=-16 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S885 N$3488 N$3490 N$3317 N$3282 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S886 N$3492 N$3494 N$3284 N$3286 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S887 N$3496 N$3498 N$3288 N$3290 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S888 N$3500 N$3504 N$3292 N$3319 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C889 N$3281 N$3283 N$3305 N$3294 "Waveguide Crossing" sch_x=-12 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C890 N$3285 N$3287 N$3296 N$3298 "Waveguide Crossing" sch_x=-12 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C891 N$3289 N$3291 N$3300 N$3315 "Waveguide Crossing" sch_x=-12 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C892 N$3293 N$3295 N$3307 N$3302 "Waveguide Crossing" sch_x=-10 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C893 N$3297 N$3299 N$3304 N$3313 "Waveguide Crossing" sch_x=-10 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C894 N$3301 N$3303 N$3309 N$3311 "Waveguide Crossing" sch_x=-8 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S833 N$3502 N$3474 N$3141 N$3106 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S834 N$3476 N$3478 N$3108 N$3110 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S835 N$3480 N$3482 N$3112 N$3114 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S836 N$3484 N$3486 N$3116 N$3143 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C837 N$3105 N$3107 N$3129 N$3118 "Waveguide Crossing" sch_x=-12 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C838 N$3109 N$3111 N$3120 N$3122 "Waveguide Crossing" sch_x=-12 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C839 N$3113 N$3115 N$3124 N$3139 "Waveguide Crossing" sch_x=-12 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C840 N$3117 N$3119 N$3131 N$3126 "Waveguide Crossing" sch_x=-10 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C841 N$3121 N$3123 N$3128 N$3137 "Waveguide Crossing" sch_x=-10 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C842 N$3125 N$3127 N$3133 N$3135 "Waveguide Crossing" sch_x=-8 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S729 N$4190 N$4130 N$2861 N$2722 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S730 N$4132 N$4134 N$2724 N$2726 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S731 N$4136 N$4138 N$2728 N$2730 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S732 N$4140 N$4142 N$2732 N$2734 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S733 N$4144 N$4146 N$2736 N$2738 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S734 N$4148 N$4150 N$2740 N$2742 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S735 N$4152 N$4154 N$2744 N$2746 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S736 N$4156 N$4158 N$2748 N$2863 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C737 N$2721 N$2723 N$2833 N$2750 "Waveguide Crossing" sch_x=-28 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C738 N$2725 N$2727 N$2752 N$2754 "Waveguide Crossing" sch_x=-28 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C739 N$2729 N$2731 N$2756 N$2758 "Waveguide Crossing" sch_x=-28 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C740 N$2733 N$2735 N$2760 N$2762 "Waveguide Crossing" sch_x=-28 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C741 N$2737 N$2739 N$2764 N$2766 "Waveguide Crossing" sch_x=-28 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C742 N$2741 N$2743 N$2768 N$2770 "Waveguide Crossing" sch_x=-28 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C743 N$2745 N$2747 N$2772 N$2859 "Waveguide Crossing" sch_x=-28 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C744 N$2749 N$2751 N$2835 N$2774 "Waveguide Crossing" sch_x=-26 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C745 N$2753 N$2755 N$2776 N$2778 "Waveguide Crossing" sch_x=-26 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C746 N$2757 N$2759 N$2780 N$2782 "Waveguide Crossing" sch_x=-26 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C747 N$2761 N$2763 N$2784 N$2786 "Waveguide Crossing" sch_x=-26 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C748 N$2765 N$2767 N$2788 N$2790 "Waveguide Crossing" sch_x=-26 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C749 N$2769 N$2771 N$2792 N$2857 "Waveguide Crossing" sch_x=-26 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C750 N$2773 N$2775 N$2837 N$2794 "Waveguide Crossing" sch_x=-24 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C751 N$2777 N$2779 N$2796 N$2798 "Waveguide Crossing" sch_x=-24 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C752 N$2781 N$2783 N$2800 N$2802 "Waveguide Crossing" sch_x=-24 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C753 N$2785 N$2787 N$2804 N$2806 "Waveguide Crossing" sch_x=-24 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C754 N$2789 N$2791 N$2808 N$2855 "Waveguide Crossing" sch_x=-24 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C755 N$2793 N$2795 N$2839 N$2810 "Waveguide Crossing" sch_x=-22 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C756 N$2797 N$2799 N$2812 N$2814 "Waveguide Crossing" sch_x=-22 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C757 N$2801 N$2803 N$2816 N$2818 "Waveguide Crossing" sch_x=-22 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C758 N$2805 N$2807 N$2820 N$2853 "Waveguide Crossing" sch_x=-22 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C759 N$2809 N$2811 N$2841 N$2822 "Waveguide Crossing" sch_x=-20 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C760 N$2813 N$2815 N$2824 N$2826 "Waveguide Crossing" sch_x=-20 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C761 N$2817 N$2819 N$2828 N$2851 "Waveguide Crossing" sch_x=-20 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C762 N$2821 N$2823 N$2843 N$2830 "Waveguide Crossing" sch_x=-18 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C763 N$2825 N$2827 N$2832 N$2849 "Waveguide Crossing" sch_x=-18 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C764 N$2829 N$2831 N$2845 N$2847 "Waveguide Crossing" sch_x=-16 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S709 N$2848 N$2850 N$2677 N$2642 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S710 N$2852 N$2854 N$2644 N$2646 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S711 N$2856 N$2858 N$2648 N$2650 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S712 N$2860 N$2864 N$2652 N$2679 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C713 N$2641 N$2643 N$2665 N$2654 "Waveguide Crossing" sch_x=-12 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C714 N$2645 N$2647 N$2656 N$2658 "Waveguide Crossing" sch_x=-12 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C715 N$2649 N$2651 N$2660 N$2675 "Waveguide Crossing" sch_x=-12 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C716 N$2653 N$2655 N$2667 N$2662 "Waveguide Crossing" sch_x=-10 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C717 N$2657 N$2659 N$2664 N$2673 "Waveguide Crossing" sch_x=-10 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C718 N$2661 N$2663 N$2669 N$2671 "Waveguide Crossing" sch_x=-8 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S657 N$2862 N$2834 N$2501 N$2466 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S658 N$2836 N$2838 N$2468 N$2470 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S659 N$2840 N$2842 N$2472 N$2474 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S660 N$2844 N$2846 N$2476 N$2503 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C661 N$2465 N$2467 N$2489 N$2478 "Waveguide Crossing" sch_x=-12 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C662 N$2469 N$2471 N$2480 N$2482 "Waveguide Crossing" sch_x=-12 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C663 N$2473 N$2475 N$2484 N$2499 "Waveguide Crossing" sch_x=-12 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C664 N$2477 N$2479 N$2491 N$2486 "Waveguide Crossing" sch_x=-10 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C665 N$2481 N$2483 N$2488 N$2497 "Waveguide Crossing" sch_x=-10 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C666 N$2485 N$2487 N$2493 N$2495 "Waveguide Crossing" sch_x=-8 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S353 N$6846 N$6722 N$1821 N$1282 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S354 N$6724 N$6726 N$1284 N$1286 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S355 N$6728 N$6730 N$1288 N$1290 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S356 N$6732 N$6734 N$1292 N$1294 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S357 N$6736 N$6738 N$1296 N$1298 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S358 N$6740 N$6742 N$1300 N$1302 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S359 N$6744 N$6746 N$1304 N$1306 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S360 N$6748 N$6750 N$1308 N$1310 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S361 N$6752 N$6754 N$1312 N$1314 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S362 N$6756 N$6758 N$1316 N$1318 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S363 N$6760 N$6762 N$1320 N$1322 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S364 N$6764 N$6766 N$1324 N$1326 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S365 N$6768 N$6770 N$1328 N$1330 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S366 N$6772 N$6774 N$1332 N$1334 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S367 N$6776 N$6778 N$1336 N$1338 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S368 N$6780 N$6782 N$1340 N$1823 MMI_switch_ideal library="Design kits/capstone" sch_x=-62 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C369 N$1281 N$1283 N$1761 N$1342 "Waveguide Crossing" sch_x=-60 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C370 N$1285 N$1287 N$1344 N$1346 "Waveguide Crossing" sch_x=-60 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C371 N$1289 N$1291 N$1348 N$1350 "Waveguide Crossing" sch_x=-60 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C372 N$1293 N$1295 N$1352 N$1354 "Waveguide Crossing" sch_x=-60 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C373 N$1297 N$1299 N$1356 N$1358 "Waveguide Crossing" sch_x=-60 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C374 N$1301 N$1303 N$1360 N$1362 "Waveguide Crossing" sch_x=-60 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C375 N$1305 N$1307 N$1364 N$1366 "Waveguide Crossing" sch_x=-60 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C376 N$1309 N$1311 N$1368 N$1370 "Waveguide Crossing" sch_x=-60 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C377 N$1313 N$1315 N$1372 N$1374 "Waveguide Crossing" sch_x=-60 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C378 N$1317 N$1319 N$1376 N$1378 "Waveguide Crossing" sch_x=-60 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C379 N$1321 N$1323 N$1380 N$1382 "Waveguide Crossing" sch_x=-60 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C380 N$1325 N$1327 N$1384 N$1386 "Waveguide Crossing" sch_x=-60 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C381 N$1329 N$1331 N$1388 N$1390 "Waveguide Crossing" sch_x=-60 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C382 N$1333 N$1335 N$1392 N$1394 "Waveguide Crossing" sch_x=-60 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C383 N$1337 N$1339 N$1396 N$1819 "Waveguide Crossing" sch_x=-60 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C384 N$1341 N$1343 N$1763 N$1398 "Waveguide Crossing" sch_x=-58 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C385 N$1345 N$1347 N$1400 N$1402 "Waveguide Crossing" sch_x=-58 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C386 N$1349 N$1351 N$1404 N$1406 "Waveguide Crossing" sch_x=-58 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C387 N$1353 N$1355 N$1408 N$1410 "Waveguide Crossing" sch_x=-58 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C388 N$1357 N$1359 N$1412 N$1414 "Waveguide Crossing" sch_x=-58 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C389 N$1361 N$1363 N$1416 N$1418 "Waveguide Crossing" sch_x=-58 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C390 N$1365 N$1367 N$1420 N$1422 "Waveguide Crossing" sch_x=-58 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C391 N$1369 N$1371 N$1424 N$1426 "Waveguide Crossing" sch_x=-58 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C392 N$1373 N$1375 N$1428 N$1430 "Waveguide Crossing" sch_x=-58 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C393 N$1377 N$1379 N$1432 N$1434 "Waveguide Crossing" sch_x=-58 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C394 N$1381 N$1383 N$1436 N$1438 "Waveguide Crossing" sch_x=-58 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C395 N$1385 N$1387 N$1440 N$1442 "Waveguide Crossing" sch_x=-58 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C396 N$1389 N$1391 N$1444 N$1446 "Waveguide Crossing" sch_x=-58 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C397 N$1393 N$1395 N$1448 N$1817 "Waveguide Crossing" sch_x=-58 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C398 N$1397 N$1399 N$1765 N$1450 "Waveguide Crossing" sch_x=-56 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C399 N$1401 N$1403 N$1452 N$1454 "Waveguide Crossing" sch_x=-56 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C400 N$1405 N$1407 N$1456 N$1458 "Waveguide Crossing" sch_x=-56 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C401 N$1409 N$1411 N$1460 N$1462 "Waveguide Crossing" sch_x=-56 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C402 N$1413 N$1415 N$1464 N$1466 "Waveguide Crossing" sch_x=-56 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C403 N$1417 N$1419 N$1468 N$1470 "Waveguide Crossing" sch_x=-56 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C404 N$1421 N$1423 N$1472 N$1474 "Waveguide Crossing" sch_x=-56 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C405 N$1425 N$1427 N$1476 N$1478 "Waveguide Crossing" sch_x=-56 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C406 N$1429 N$1431 N$1480 N$1482 "Waveguide Crossing" sch_x=-56 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C407 N$1433 N$1435 N$1484 N$1486 "Waveguide Crossing" sch_x=-56 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C408 N$1437 N$1439 N$1488 N$1490 "Waveguide Crossing" sch_x=-56 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C409 N$1441 N$1443 N$1492 N$1494 "Waveguide Crossing" sch_x=-56 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C410 N$1445 N$1447 N$1496 N$1815 "Waveguide Crossing" sch_x=-56 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C411 N$1449 N$1451 N$1767 N$1498 "Waveguide Crossing" sch_x=-54 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C412 N$1453 N$1455 N$1500 N$1502 "Waveguide Crossing" sch_x=-54 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C413 N$1457 N$1459 N$1504 N$1506 "Waveguide Crossing" sch_x=-54 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C414 N$1461 N$1463 N$1508 N$1510 "Waveguide Crossing" sch_x=-54 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C415 N$1465 N$1467 N$1512 N$1514 "Waveguide Crossing" sch_x=-54 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C416 N$1469 N$1471 N$1516 N$1518 "Waveguide Crossing" sch_x=-54 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C417 N$1473 N$1475 N$1520 N$1522 "Waveguide Crossing" sch_x=-54 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C418 N$1477 N$1479 N$1524 N$1526 "Waveguide Crossing" sch_x=-54 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C419 N$1481 N$1483 N$1528 N$1530 "Waveguide Crossing" sch_x=-54 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C420 N$1485 N$1487 N$1532 N$1534 "Waveguide Crossing" sch_x=-54 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C421 N$1489 N$1491 N$1536 N$1538 "Waveguide Crossing" sch_x=-54 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C422 N$1493 N$1495 N$1540 N$1813 "Waveguide Crossing" sch_x=-54 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C423 N$1497 N$1499 N$1769 N$1542 "Waveguide Crossing" sch_x=-52 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C424 N$1501 N$1503 N$1544 N$1546 "Waveguide Crossing" sch_x=-52 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C425 N$1505 N$1507 N$1548 N$1550 "Waveguide Crossing" sch_x=-52 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C426 N$1509 N$1511 N$1552 N$1554 "Waveguide Crossing" sch_x=-52 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C427 N$1513 N$1515 N$1556 N$1558 "Waveguide Crossing" sch_x=-52 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C428 N$1517 N$1519 N$1560 N$1562 "Waveguide Crossing" sch_x=-52 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C429 N$1521 N$1523 N$1564 N$1566 "Waveguide Crossing" sch_x=-52 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C430 N$1525 N$1527 N$1568 N$1570 "Waveguide Crossing" sch_x=-52 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C431 N$1529 N$1531 N$1572 N$1574 "Waveguide Crossing" sch_x=-52 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C432 N$1533 N$1535 N$1576 N$1578 "Waveguide Crossing" sch_x=-52 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C433 N$1537 N$1539 N$1580 N$1811 "Waveguide Crossing" sch_x=-52 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C434 N$1541 N$1543 N$1771 N$1582 "Waveguide Crossing" sch_x=-50 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C435 N$1545 N$1547 N$1584 N$1586 "Waveguide Crossing" sch_x=-50 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C436 N$1549 N$1551 N$1588 N$1590 "Waveguide Crossing" sch_x=-50 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C437 N$1553 N$1555 N$1592 N$1594 "Waveguide Crossing" sch_x=-50 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C438 N$1557 N$1559 N$1596 N$1598 "Waveguide Crossing" sch_x=-50 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C439 N$1561 N$1563 N$1600 N$1602 "Waveguide Crossing" sch_x=-50 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C440 N$1565 N$1567 N$1604 N$1606 "Waveguide Crossing" sch_x=-50 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C441 N$1569 N$1571 N$1608 N$1610 "Waveguide Crossing" sch_x=-50 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C442 N$1573 N$1575 N$1612 N$1614 "Waveguide Crossing" sch_x=-50 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C443 N$1577 N$1579 N$1616 N$1809 "Waveguide Crossing" sch_x=-50 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C444 N$1581 N$1583 N$1773 N$1618 "Waveguide Crossing" sch_x=-48 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C445 N$1585 N$1587 N$1620 N$1622 "Waveguide Crossing" sch_x=-48 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C446 N$1589 N$1591 N$1624 N$1626 "Waveguide Crossing" sch_x=-48 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C447 N$1593 N$1595 N$1628 N$1630 "Waveguide Crossing" sch_x=-48 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C448 N$1597 N$1599 N$1632 N$1634 "Waveguide Crossing" sch_x=-48 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C449 N$1601 N$1603 N$1636 N$1638 "Waveguide Crossing" sch_x=-48 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C450 N$1605 N$1607 N$1640 N$1642 "Waveguide Crossing" sch_x=-48 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C451 N$1609 N$1611 N$1644 N$1646 "Waveguide Crossing" sch_x=-48 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C452 N$1613 N$1615 N$1648 N$1807 "Waveguide Crossing" sch_x=-48 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C453 N$1617 N$1619 N$1775 N$1650 "Waveguide Crossing" sch_x=-46 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C454 N$1621 N$1623 N$1652 N$1654 "Waveguide Crossing" sch_x=-46 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C455 N$1625 N$1627 N$1656 N$1658 "Waveguide Crossing" sch_x=-46 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C456 N$1629 N$1631 N$1660 N$1662 "Waveguide Crossing" sch_x=-46 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C457 N$1633 N$1635 N$1664 N$1666 "Waveguide Crossing" sch_x=-46 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C458 N$1637 N$1639 N$1668 N$1670 "Waveguide Crossing" sch_x=-46 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C459 N$1641 N$1643 N$1672 N$1674 "Waveguide Crossing" sch_x=-46 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C460 N$1645 N$1647 N$1676 N$1805 "Waveguide Crossing" sch_x=-46 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C461 N$1649 N$1651 N$1777 N$1678 "Waveguide Crossing" sch_x=-44 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C462 N$1653 N$1655 N$1680 N$1682 "Waveguide Crossing" sch_x=-44 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C463 N$1657 N$1659 N$1684 N$1686 "Waveguide Crossing" sch_x=-44 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C464 N$1661 N$1663 N$1688 N$1690 "Waveguide Crossing" sch_x=-44 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C465 N$1665 N$1667 N$1692 N$1694 "Waveguide Crossing" sch_x=-44 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C466 N$1669 N$1671 N$1696 N$1698 "Waveguide Crossing" sch_x=-44 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C467 N$1673 N$1675 N$1700 N$1803 "Waveguide Crossing" sch_x=-44 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C468 N$1677 N$1679 N$1779 N$1702 "Waveguide Crossing" sch_x=-42 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C469 N$1681 N$1683 N$1704 N$1706 "Waveguide Crossing" sch_x=-42 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C470 N$1685 N$1687 N$1708 N$1710 "Waveguide Crossing" sch_x=-42 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C471 N$1689 N$1691 N$1712 N$1714 "Waveguide Crossing" sch_x=-42 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C472 N$1693 N$1695 N$1716 N$1718 "Waveguide Crossing" sch_x=-42 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C473 N$1697 N$1699 N$1720 N$1801 "Waveguide Crossing" sch_x=-42 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C474 N$1701 N$1703 N$1781 N$1722 "Waveguide Crossing" sch_x=-40 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C475 N$1705 N$1707 N$1724 N$1726 "Waveguide Crossing" sch_x=-40 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C476 N$1709 N$1711 N$1728 N$1730 "Waveguide Crossing" sch_x=-40 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C477 N$1713 N$1715 N$1732 N$1734 "Waveguide Crossing" sch_x=-40 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C478 N$1717 N$1719 N$1736 N$1799 "Waveguide Crossing" sch_x=-40 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C479 N$1721 N$1723 N$1783 N$1738 "Waveguide Crossing" sch_x=-38 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C480 N$1725 N$1727 N$1740 N$1742 "Waveguide Crossing" sch_x=-38 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C481 N$1729 N$1731 N$1744 N$1746 "Waveguide Crossing" sch_x=-38 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C482 N$1733 N$1735 N$1748 N$1797 "Waveguide Crossing" sch_x=-38 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C483 N$1737 N$1739 N$1785 N$1750 "Waveguide Crossing" sch_x=-36 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C484 N$1741 N$1743 N$1752 N$1754 "Waveguide Crossing" sch_x=-36 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C485 N$1745 N$1747 N$1756 N$1795 "Waveguide Crossing" sch_x=-36 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C486 N$1749 N$1751 N$1787 N$1758 "Waveguide Crossing" sch_x=-34 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C487 N$1753 N$1755 N$1760 N$1793 "Waveguide Crossing" sch_x=-34 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C488 N$1757 N$1759 N$1789 N$1791 "Waveguide Crossing" sch_x=-32 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S281 N$1792 N$1794 N$1133 N$994 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S282 N$1796 N$1798 N$996 N$998 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S283 N$1800 N$1802 N$1000 N$1002 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S284 N$1804 N$1806 N$1004 N$1006 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S285 N$1808 N$1810 N$1008 N$1010 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S286 N$1812 N$1814 N$1012 N$1014 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S287 N$1816 N$1818 N$1016 N$1018 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S288 N$1820 N$1824 N$1020 N$1135 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C289 N$993 N$995 N$1105 N$1022 "Waveguide Crossing" sch_x=-28 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C290 N$997 N$999 N$1024 N$1026 "Waveguide Crossing" sch_x=-28 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C291 N$1001 N$1003 N$1028 N$1030 "Waveguide Crossing" sch_x=-28 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C292 N$1005 N$1007 N$1032 N$1034 "Waveguide Crossing" sch_x=-28 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C293 N$1009 N$1011 N$1036 N$1038 "Waveguide Crossing" sch_x=-28 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C294 N$1013 N$1015 N$1040 N$1042 "Waveguide Crossing" sch_x=-28 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C295 N$1017 N$1019 N$1044 N$1131 "Waveguide Crossing" sch_x=-28 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C296 N$1021 N$1023 N$1107 N$1046 "Waveguide Crossing" sch_x=-26 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C297 N$1025 N$1027 N$1048 N$1050 "Waveguide Crossing" sch_x=-26 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C298 N$1029 N$1031 N$1052 N$1054 "Waveguide Crossing" sch_x=-26 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C299 N$1033 N$1035 N$1056 N$1058 "Waveguide Crossing" sch_x=-26 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C300 N$1037 N$1039 N$1060 N$1062 "Waveguide Crossing" sch_x=-26 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C301 N$1041 N$1043 N$1064 N$1129 "Waveguide Crossing" sch_x=-26 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C302 N$1045 N$1047 N$1109 N$1066 "Waveguide Crossing" sch_x=-24 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C303 N$1049 N$1051 N$1068 N$1070 "Waveguide Crossing" sch_x=-24 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C304 N$1053 N$1055 N$1072 N$1074 "Waveguide Crossing" sch_x=-24 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C305 N$1057 N$1059 N$1076 N$1078 "Waveguide Crossing" sch_x=-24 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C306 N$1061 N$1063 N$1080 N$1127 "Waveguide Crossing" sch_x=-24 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C307 N$1065 N$1067 N$1111 N$1082 "Waveguide Crossing" sch_x=-22 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C308 N$1069 N$1071 N$1084 N$1086 "Waveguide Crossing" sch_x=-22 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C309 N$1073 N$1075 N$1088 N$1090 "Waveguide Crossing" sch_x=-22 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C310 N$1077 N$1079 N$1092 N$1125 "Waveguide Crossing" sch_x=-22 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C311 N$1081 N$1083 N$1113 N$1094 "Waveguide Crossing" sch_x=-20 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C312 N$1085 N$1087 N$1096 N$1098 "Waveguide Crossing" sch_x=-20 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C313 N$1089 N$1091 N$1100 N$1123 "Waveguide Crossing" sch_x=-20 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C314 N$1093 N$1095 N$1115 N$1102 "Waveguide Crossing" sch_x=-18 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C315 N$1097 N$1099 N$1104 N$1121 "Waveguide Crossing" sch_x=-18 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C316 N$1101 N$1103 N$1117 N$1119 "Waveguide Crossing" sch_x=-16 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S261 N$1120 N$1122 N$949 N$914 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S262 N$1124 N$1126 N$916 N$918 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S263 N$1128 N$1130 N$920 N$922 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S264 N$1132 N$1136 N$924 N$951 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C265 N$913 N$915 N$937 N$926 "Waveguide Crossing" sch_x=-12 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C266 N$917 N$919 N$928 N$930 "Waveguide Crossing" sch_x=-12 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C267 N$921 N$923 N$932 N$947 "Waveguide Crossing" sch_x=-12 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C268 N$925 N$927 N$939 N$934 "Waveguide Crossing" sch_x=-10 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C269 N$929 N$931 N$936 N$945 "Waveguide Crossing" sch_x=-10 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C270 N$933 N$935 N$941 N$943 "Waveguide Crossing" sch_x=-8 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S209 N$1134 N$1106 N$773 N$738 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S210 N$1108 N$1110 N$740 N$742 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S211 N$1112 N$1114 N$744 N$746 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S212 N$1116 N$1118 N$748 N$775 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C213 N$737 N$739 N$761 N$750 "Waveguide Crossing" sch_x=-12 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C214 N$741 N$743 N$752 N$754 "Waveguide Crossing" sch_x=-12 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C215 N$745 N$747 N$756 N$771 "Waveguide Crossing" sch_x=-12 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C216 N$749 N$751 N$763 N$758 "Waveguide Crossing" sch_x=-10 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C217 N$753 N$755 N$760 N$769 "Waveguide Crossing" sch_x=-10 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C218 N$757 N$759 N$765 N$767 "Waveguide Crossing" sch_x=-8 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S105 N$1822 N$1762 N$493 N$354 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S106 N$1764 N$1766 N$356 N$358 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S107 N$1768 N$1770 N$360 N$362 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S108 N$1772 N$1774 N$364 N$366 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S109 N$1776 N$1778 N$368 N$370 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S110 N$1780 N$1782 N$372 N$374 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S111 N$1784 N$1786 N$376 N$378 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S112 N$1788 N$1790 N$380 N$495 MMI_switch_ideal library="Design kits/capstone" sch_x=-30 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C113 N$353 N$355 N$465 N$382 "Waveguide Crossing" sch_x=-28 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C114 N$357 N$359 N$384 N$386 "Waveguide Crossing" sch_x=-28 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C115 N$361 N$363 N$388 N$390 "Waveguide Crossing" sch_x=-28 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C116 N$365 N$367 N$392 N$394 "Waveguide Crossing" sch_x=-28 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C117 N$369 N$371 N$396 N$398 "Waveguide Crossing" sch_x=-28 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C118 N$373 N$375 N$400 N$402 "Waveguide Crossing" sch_x=-28 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C119 N$377 N$379 N$404 N$491 "Waveguide Crossing" sch_x=-28 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C120 N$381 N$383 N$467 N$406 "Waveguide Crossing" sch_x=-26 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C121 N$385 N$387 N$408 N$410 "Waveguide Crossing" sch_x=-26 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C122 N$389 N$391 N$412 N$414 "Waveguide Crossing" sch_x=-26 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C123 N$393 N$395 N$416 N$418 "Waveguide Crossing" sch_x=-26 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C124 N$397 N$399 N$420 N$422 "Waveguide Crossing" sch_x=-26 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C125 N$401 N$403 N$424 N$489 "Waveguide Crossing" sch_x=-26 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C126 N$405 N$407 N$469 N$426 "Waveguide Crossing" sch_x=-24 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C127 N$409 N$411 N$428 N$430 "Waveguide Crossing" sch_x=-24 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C128 N$413 N$415 N$432 N$434 "Waveguide Crossing" sch_x=-24 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C129 N$417 N$419 N$436 N$438 "Waveguide Crossing" sch_x=-24 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C130 N$421 N$423 N$440 N$487 "Waveguide Crossing" sch_x=-24 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C131 N$425 N$427 N$471 N$442 "Waveguide Crossing" sch_x=-22 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C132 N$429 N$431 N$444 N$446 "Waveguide Crossing" sch_x=-22 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C133 N$433 N$435 N$448 N$450 "Waveguide Crossing" sch_x=-22 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C134 N$437 N$439 N$452 N$485 "Waveguide Crossing" sch_x=-22 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C135 N$441 N$443 N$473 N$454 "Waveguide Crossing" sch_x=-20 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C136 N$445 N$447 N$456 N$458 "Waveguide Crossing" sch_x=-20 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C137 N$449 N$451 N$460 N$483 "Waveguide Crossing" sch_x=-20 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C138 N$453 N$455 N$475 N$462 "Waveguide Crossing" sch_x=-18 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C139 N$457 N$459 N$464 N$481 "Waveguide Crossing" sch_x=-18 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C140 N$461 N$463 N$477 N$479 "Waveguide Crossing" sch_x=-16 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S85 N$480 N$482 N$309 N$274 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S86 N$484 N$486 N$276 N$278 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S87 N$488 N$490 N$280 N$282 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S88 N$492 N$496 N$284 N$311 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C89 N$273 N$275 N$297 N$286 "Waveguide Crossing" sch_x=-12 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C90 N$277 N$279 N$288 N$290 "Waveguide Crossing" sch_x=-12 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C91 N$281 N$283 N$292 N$307 "Waveguide Crossing" sch_x=-12 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C92 N$285 N$287 N$299 N$294 "Waveguide Crossing" sch_x=-10 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C93 N$289 N$291 N$296 N$305 "Waveguide Crossing" sch_x=-10 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C94 N$293 N$295 N$301 N$303 "Waveguide Crossing" sch_x=-8 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S33 N$494 N$466 N$133 N$98 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S34 N$468 N$470 N$100 N$102 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S35 N$472 N$474 N$104 N$106 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S36 N$476 N$478 N$108 N$135 MMI_switch_ideal library="Design kits/capstone" sch_x=-14 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C37 N$97 N$99 N$121 N$110 "Waveguide Crossing" sch_x=-12 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C38 N$101 N$103 N$112 N$114 "Waveguide Crossing" sch_x=-12 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C39 N$105 N$107 N$116 N$131 "Waveguide Crossing" sch_x=-12 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C40 N$109 N$111 N$123 N$118 "Waveguide Crossing" sch_x=-10 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C41 N$113 N$115 N$120 N$129 "Waveguide Crossing" sch_x=-10 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C42 N$117 N$119 N$125 N$127 "Waveguide Crossing" sch_x=-8 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1 N$134 N$122 N$1 N$3 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2 N$124 N$126 N$5 N$11 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3 N$9025 N$2 N$13 N$15 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4 N$8 N$9026 N$17 N$23 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S5 N$9027 N$10 N$25 N$27 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6 N$12 N$9028 N$29 N$35 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S7 N$14 N$22 N$37 N$9029 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S8 N$20 N$24 N$9030 N$39 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S9 N$26 N$34 N$41 N$9031 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S10 N$32 N$36 N$9032 N$47 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S11 N$38 N$46 N$174 N$162 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S12 N$44 N$48 N$164 N$166 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C13 N$4 N$6 N$7 N$9 "Waveguide Crossing" sch_x=-4 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C14 N$16 N$18 N$21 N$19 "Waveguide Crossing" sch_x=0 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C15 N$28 N$30 N$33 N$31 "Waveguide Crossing" sch_x=0 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C16 N$40 N$42 N$45 N$43 "Waveguide Crossing" sch_x=4 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S17 N$128 N$130 N$49 N$51 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S18 N$132 N$136 N$53 N$59 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S19 N$9033 N$50 N$61 N$63 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S20 N$56 N$9034 N$65 N$71 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S21 N$9035 N$58 N$73 N$75 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S22 N$60 N$9036 N$77 N$83 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S23 N$62 N$70 N$85 N$9037 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S24 N$68 N$72 N$9038 N$87 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S25 N$74 N$82 N$89 N$9039 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S26 N$80 N$84 N$9040 N$95 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S27 N$86 N$94 N$168 N$170 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S28 N$92 N$96 N$172 N$176 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C29 N$52 N$54 N$55 N$57 "Waveguide Crossing" sch_x=-4 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C30 N$64 N$66 N$69 N$67 "Waveguide Crossing" sch_x=0 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C31 N$76 N$78 N$81 N$79 "Waveguide Crossing" sch_x=0 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C32 N$88 N$90 N$93 N$91 "Waveguide Crossing" sch_x=4 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C47 N$161 N$150 N$137 N$139 "Waveguide Crossing" sch_x=12 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C48 N$152 N$154 N$141 N$143 "Waveguide Crossing" sch_x=12 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C49 N$156 N$171 N$145 N$147 "Waveguide Crossing" sch_x=12 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C50 N$163 N$158 N$149 N$151 "Waveguide Crossing" sch_x=10 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C51 N$160 N$169 N$153 N$155 "Waveguide Crossing" sch_x=10 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C52 N$165 N$167 N$157 N$159 "Waveguide Crossing" sch_x=8 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S43 N$173 N$138 N$638 N$610 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S44 N$140 N$142 N$612 N$614 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S45 N$144 N$146 N$616 N$618 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S46 N$148 N$175 N$620 N$622 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S53 N$310 N$298 N$177 N$179 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S54 N$300 N$302 N$181 N$187 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S55 N$9041 N$178 N$189 N$191 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S56 N$184 N$9042 N$193 N$199 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S57 N$9043 N$186 N$201 N$203 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S58 N$188 N$9044 N$205 N$211 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S59 N$190 N$198 N$213 N$9045 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S60 N$196 N$200 N$9046 N$215 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S61 N$202 N$210 N$217 N$9047 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S62 N$208 N$212 N$9048 N$223 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S63 N$214 N$222 N$350 N$338 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S64 N$220 N$224 N$340 N$342 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C65 N$180 N$182 N$183 N$185 "Waveguide Crossing" sch_x=-4 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C66 N$192 N$194 N$197 N$195 "Waveguide Crossing" sch_x=0 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C67 N$204 N$206 N$209 N$207 "Waveguide Crossing" sch_x=0 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C68 N$216 N$218 N$221 N$219 "Waveguide Crossing" sch_x=4 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S69 N$304 N$306 N$225 N$227 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S70 N$308 N$312 N$229 N$235 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S71 N$9049 N$226 N$237 N$239 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S72 N$232 N$9050 N$241 N$247 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S73 N$9051 N$234 N$249 N$251 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S74 N$236 N$9052 N$253 N$259 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S75 N$238 N$246 N$261 N$9053 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S76 N$244 N$248 N$9054 N$263 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S77 N$250 N$258 N$265 N$9055 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S78 N$256 N$260 N$9056 N$271 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S79 N$262 N$270 N$344 N$346 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S80 N$268 N$272 N$348 N$352 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C81 N$228 N$230 N$231 N$233 "Waveguide Crossing" sch_x=-4 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C82 N$240 N$242 N$245 N$243 "Waveguide Crossing" sch_x=0 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C83 N$252 N$254 N$257 N$255 "Waveguide Crossing" sch_x=0 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C84 N$264 N$266 N$269 N$267 "Waveguide Crossing" sch_x=4 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C99 N$337 N$326 N$313 N$315 "Waveguide Crossing" sch_x=12 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C100 N$328 N$330 N$317 N$319 "Waveguide Crossing" sch_x=12 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C101 N$332 N$347 N$321 N$323 "Waveguide Crossing" sch_x=12 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C102 N$339 N$334 N$325 N$327 "Waveguide Crossing" sch_x=10 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C103 N$336 N$345 N$329 N$331 "Waveguide Crossing" sch_x=10 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C104 N$341 N$343 N$333 N$335 "Waveguide Crossing" sch_x=8 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S95 N$349 N$314 N$624 N$626 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S96 N$316 N$318 N$628 N$630 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S97 N$320 N$322 N$632 N$634 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S98 N$324 N$351 N$636 N$640 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C149 N$609 N$526 N$497 N$499 "Waveguide Crossing" sch_x=28 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C150 N$528 N$530 N$501 N$503 "Waveguide Crossing" sch_x=28 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C151 N$532 N$534 N$505 N$507 "Waveguide Crossing" sch_x=28 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C152 N$536 N$538 N$509 N$511 "Waveguide Crossing" sch_x=28 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C153 N$540 N$542 N$513 N$515 "Waveguide Crossing" sch_x=28 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C154 N$544 N$546 N$517 N$519 "Waveguide Crossing" sch_x=28 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C155 N$548 N$635 N$521 N$523 "Waveguide Crossing" sch_x=28 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C156 N$611 N$550 N$525 N$527 "Waveguide Crossing" sch_x=26 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C157 N$552 N$554 N$529 N$531 "Waveguide Crossing" sch_x=26 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C158 N$556 N$558 N$533 N$535 "Waveguide Crossing" sch_x=26 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C159 N$560 N$562 N$537 N$539 "Waveguide Crossing" sch_x=26 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C160 N$564 N$566 N$541 N$543 "Waveguide Crossing" sch_x=26 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C161 N$568 N$633 N$545 N$547 "Waveguide Crossing" sch_x=26 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C162 N$613 N$570 N$549 N$551 "Waveguide Crossing" sch_x=24 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C163 N$572 N$574 N$553 N$555 "Waveguide Crossing" sch_x=24 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C164 N$576 N$578 N$557 N$559 "Waveguide Crossing" sch_x=24 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C165 N$580 N$582 N$561 N$563 "Waveguide Crossing" sch_x=24 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C166 N$584 N$631 N$565 N$567 "Waveguide Crossing" sch_x=24 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C167 N$615 N$586 N$569 N$571 "Waveguide Crossing" sch_x=22 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C168 N$588 N$590 N$573 N$575 "Waveguide Crossing" sch_x=22 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C169 N$592 N$594 N$577 N$579 "Waveguide Crossing" sch_x=22 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C170 N$596 N$629 N$581 N$583 "Waveguide Crossing" sch_x=22 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C171 N$617 N$598 N$585 N$587 "Waveguide Crossing" sch_x=20 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C172 N$600 N$602 N$589 N$591 "Waveguide Crossing" sch_x=20 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C173 N$604 N$627 N$593 N$595 "Waveguide Crossing" sch_x=20 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C174 N$619 N$606 N$597 N$599 "Waveguide Crossing" sch_x=18 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C175 N$608 N$625 N$601 N$603 "Waveguide Crossing" sch_x=18 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C176 N$621 N$623 N$605 N$607 "Waveguide Crossing" sch_x=16 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S141 N$637 N$498 N$2366 N$2306 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S142 N$500 N$502 N$2308 N$2310 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S143 N$504 N$506 N$2312 N$2314 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S144 N$508 N$510 N$2316 N$2318 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S145 N$512 N$514 N$2320 N$2322 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S146 N$516 N$518 N$2324 N$2326 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S147 N$520 N$522 N$2328 N$2330 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S148 N$524 N$639 N$2332 N$2334 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S177 N$774 N$762 N$641 N$643 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S178 N$764 N$766 N$645 N$651 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S179 N$9057 N$642 N$653 N$655 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S180 N$648 N$9058 N$657 N$663 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S181 N$9059 N$650 N$665 N$667 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S182 N$652 N$9060 N$669 N$675 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S183 N$654 N$662 N$677 N$9061 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S184 N$660 N$664 N$9062 N$679 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S185 N$666 N$674 N$681 N$9063 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S186 N$672 N$676 N$9064 N$687 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S187 N$678 N$686 N$814 N$802 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S188 N$684 N$688 N$804 N$806 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C189 N$644 N$646 N$647 N$649 "Waveguide Crossing" sch_x=-4 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C190 N$656 N$658 N$661 N$659 "Waveguide Crossing" sch_x=0 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C191 N$668 N$670 N$673 N$671 "Waveguide Crossing" sch_x=0 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C192 N$680 N$682 N$685 N$683 "Waveguide Crossing" sch_x=4 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S193 N$768 N$770 N$689 N$691 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S194 N$772 N$776 N$693 N$699 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S195 N$9065 N$690 N$701 N$703 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S196 N$696 N$9066 N$705 N$711 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S197 N$9067 N$698 N$713 N$715 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S198 N$700 N$9068 N$717 N$723 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S199 N$702 N$710 N$725 N$9069 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S200 N$708 N$712 N$9070 N$727 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S201 N$714 N$722 N$729 N$9071 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S202 N$720 N$724 N$9072 N$735 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S203 N$726 N$734 N$808 N$810 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S204 N$732 N$736 N$812 N$816 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C205 N$692 N$694 N$695 N$697 "Waveguide Crossing" sch_x=-4 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C206 N$704 N$706 N$709 N$707 "Waveguide Crossing" sch_x=0 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C207 N$716 N$718 N$721 N$719 "Waveguide Crossing" sch_x=0 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C208 N$728 N$730 N$733 N$731 "Waveguide Crossing" sch_x=4 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C223 N$801 N$790 N$777 N$779 "Waveguide Crossing" sch_x=12 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C224 N$792 N$794 N$781 N$783 "Waveguide Crossing" sch_x=12 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C225 N$796 N$811 N$785 N$787 "Waveguide Crossing" sch_x=12 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C226 N$803 N$798 N$789 N$791 "Waveguide Crossing" sch_x=10 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C227 N$800 N$809 N$793 N$795 "Waveguide Crossing" sch_x=10 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C228 N$805 N$807 N$797 N$799 "Waveguide Crossing" sch_x=8 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S219 N$813 N$778 N$1278 N$1250 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S220 N$780 N$782 N$1252 N$1254 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S221 N$784 N$786 N$1256 N$1258 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S222 N$788 N$815 N$1260 N$1262 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S229 N$950 N$938 N$817 N$819 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S230 N$940 N$942 N$821 N$827 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S231 N$9073 N$818 N$829 N$831 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S232 N$824 N$9074 N$833 N$839 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S233 N$9075 N$826 N$841 N$843 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S234 N$828 N$9076 N$845 N$851 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S235 N$830 N$838 N$853 N$9077 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S236 N$836 N$840 N$9078 N$855 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S237 N$842 N$850 N$857 N$9079 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S238 N$848 N$852 N$9080 N$863 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S239 N$854 N$862 N$990 N$978 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S240 N$860 N$864 N$980 N$982 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C241 N$820 N$822 N$823 N$825 "Waveguide Crossing" sch_x=-4 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C242 N$832 N$834 N$837 N$835 "Waveguide Crossing" sch_x=0 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C243 N$844 N$846 N$849 N$847 "Waveguide Crossing" sch_x=0 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C244 N$856 N$858 N$861 N$859 "Waveguide Crossing" sch_x=4 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S245 N$944 N$946 N$865 N$867 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S246 N$948 N$952 N$869 N$875 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S247 N$9081 N$866 N$877 N$879 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S248 N$872 N$9082 N$881 N$887 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S249 N$9083 N$874 N$889 N$891 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S250 N$876 N$9084 N$893 N$899 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S251 N$878 N$886 N$901 N$9085 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S252 N$884 N$888 N$9086 N$903 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S253 N$890 N$898 N$905 N$9087 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S254 N$896 N$900 N$9088 N$911 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S255 N$902 N$910 N$984 N$986 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S256 N$908 N$912 N$988 N$992 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C257 N$868 N$870 N$871 N$873 "Waveguide Crossing" sch_x=-4 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C258 N$880 N$882 N$885 N$883 "Waveguide Crossing" sch_x=0 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C259 N$892 N$894 N$897 N$895 "Waveguide Crossing" sch_x=0 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C260 N$904 N$906 N$909 N$907 "Waveguide Crossing" sch_x=4 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C275 N$977 N$966 N$953 N$955 "Waveguide Crossing" sch_x=12 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C276 N$968 N$970 N$957 N$959 "Waveguide Crossing" sch_x=12 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C277 N$972 N$987 N$961 N$963 "Waveguide Crossing" sch_x=12 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C278 N$979 N$974 N$965 N$967 "Waveguide Crossing" sch_x=10 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C279 N$976 N$985 N$969 N$971 "Waveguide Crossing" sch_x=10 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C280 N$981 N$983 N$973 N$975 "Waveguide Crossing" sch_x=8 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S271 N$989 N$954 N$1264 N$1266 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S272 N$956 N$958 N$1268 N$1270 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S273 N$960 N$962 N$1272 N$1274 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S274 N$964 N$991 N$1276 N$1280 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C325 N$1249 N$1166 N$1137 N$1139 "Waveguide Crossing" sch_x=28 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C326 N$1168 N$1170 N$1141 N$1143 "Waveguide Crossing" sch_x=28 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C327 N$1172 N$1174 N$1145 N$1147 "Waveguide Crossing" sch_x=28 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C328 N$1176 N$1178 N$1149 N$1151 "Waveguide Crossing" sch_x=28 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C329 N$1180 N$1182 N$1153 N$1155 "Waveguide Crossing" sch_x=28 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C330 N$1184 N$1186 N$1157 N$1159 "Waveguide Crossing" sch_x=28 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C331 N$1188 N$1275 N$1161 N$1163 "Waveguide Crossing" sch_x=28 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C332 N$1251 N$1190 N$1165 N$1167 "Waveguide Crossing" sch_x=26 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C333 N$1192 N$1194 N$1169 N$1171 "Waveguide Crossing" sch_x=26 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C334 N$1196 N$1198 N$1173 N$1175 "Waveguide Crossing" sch_x=26 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C335 N$1200 N$1202 N$1177 N$1179 "Waveguide Crossing" sch_x=26 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C336 N$1204 N$1206 N$1181 N$1183 "Waveguide Crossing" sch_x=26 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C337 N$1208 N$1273 N$1185 N$1187 "Waveguide Crossing" sch_x=26 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C338 N$1253 N$1210 N$1189 N$1191 "Waveguide Crossing" sch_x=24 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C339 N$1212 N$1214 N$1193 N$1195 "Waveguide Crossing" sch_x=24 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C340 N$1216 N$1218 N$1197 N$1199 "Waveguide Crossing" sch_x=24 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C341 N$1220 N$1222 N$1201 N$1203 "Waveguide Crossing" sch_x=24 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C342 N$1224 N$1271 N$1205 N$1207 "Waveguide Crossing" sch_x=24 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C343 N$1255 N$1226 N$1209 N$1211 "Waveguide Crossing" sch_x=22 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C344 N$1228 N$1230 N$1213 N$1215 "Waveguide Crossing" sch_x=22 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C345 N$1232 N$1234 N$1217 N$1219 "Waveguide Crossing" sch_x=22 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C346 N$1236 N$1269 N$1221 N$1223 "Waveguide Crossing" sch_x=22 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C347 N$1257 N$1238 N$1225 N$1227 "Waveguide Crossing" sch_x=20 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C348 N$1240 N$1242 N$1229 N$1231 "Waveguide Crossing" sch_x=20 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C349 N$1244 N$1267 N$1233 N$1235 "Waveguide Crossing" sch_x=20 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C350 N$1259 N$1246 N$1237 N$1239 "Waveguide Crossing" sch_x=18 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C351 N$1248 N$1265 N$1241 N$1243 "Waveguide Crossing" sch_x=18 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C352 N$1261 N$1263 N$1245 N$1247 "Waveguide Crossing" sch_x=16 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S317 N$1277 N$1138 N$2336 N$2338 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S318 N$1140 N$1142 N$2340 N$2342 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S319 N$1144 N$1146 N$2344 N$2346 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S320 N$1148 N$1150 N$2348 N$2350 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S321 N$1152 N$1154 N$2352 N$2354 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S322 N$1156 N$1158 N$2356 N$2358 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S323 N$1160 N$1162 N$2360 N$2362 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S324 N$1164 N$1279 N$2364 N$2368 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C505 N$2305 N$1886 N$1825 N$1827 "Waveguide Crossing" sch_x=60 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C506 N$1888 N$1890 N$1829 N$1831 "Waveguide Crossing" sch_x=60 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C507 N$1892 N$1894 N$1833 N$1835 "Waveguide Crossing" sch_x=60 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C508 N$1896 N$1898 N$1837 N$1839 "Waveguide Crossing" sch_x=60 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C509 N$1900 N$1902 N$1841 N$1843 "Waveguide Crossing" sch_x=60 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C510 N$1904 N$1906 N$1845 N$1847 "Waveguide Crossing" sch_x=60 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C511 N$1908 N$1910 N$1849 N$1851 "Waveguide Crossing" sch_x=60 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C512 N$1912 N$1914 N$1853 N$1855 "Waveguide Crossing" sch_x=60 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C513 N$1916 N$1918 N$1857 N$1859 "Waveguide Crossing" sch_x=60 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C514 N$1920 N$1922 N$1861 N$1863 "Waveguide Crossing" sch_x=60 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C515 N$1924 N$1926 N$1865 N$1867 "Waveguide Crossing" sch_x=60 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C516 N$1928 N$1930 N$1869 N$1871 "Waveguide Crossing" sch_x=60 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C517 N$1932 N$1934 N$1873 N$1875 "Waveguide Crossing" sch_x=60 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C518 N$1936 N$1938 N$1877 N$1879 "Waveguide Crossing" sch_x=60 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C519 N$1940 N$2363 N$1881 N$1883 "Waveguide Crossing" sch_x=60 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C520 N$2307 N$1942 N$1885 N$1887 "Waveguide Crossing" sch_x=58 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C521 N$1944 N$1946 N$1889 N$1891 "Waveguide Crossing" sch_x=58 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C522 N$1948 N$1950 N$1893 N$1895 "Waveguide Crossing" sch_x=58 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C523 N$1952 N$1954 N$1897 N$1899 "Waveguide Crossing" sch_x=58 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C524 N$1956 N$1958 N$1901 N$1903 "Waveguide Crossing" sch_x=58 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C525 N$1960 N$1962 N$1905 N$1907 "Waveguide Crossing" sch_x=58 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C526 N$1964 N$1966 N$1909 N$1911 "Waveguide Crossing" sch_x=58 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C527 N$1968 N$1970 N$1913 N$1915 "Waveguide Crossing" sch_x=58 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C528 N$1972 N$1974 N$1917 N$1919 "Waveguide Crossing" sch_x=58 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C529 N$1976 N$1978 N$1921 N$1923 "Waveguide Crossing" sch_x=58 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C530 N$1980 N$1982 N$1925 N$1927 "Waveguide Crossing" sch_x=58 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C531 N$1984 N$1986 N$1929 N$1931 "Waveguide Crossing" sch_x=58 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C532 N$1988 N$1990 N$1933 N$1935 "Waveguide Crossing" sch_x=58 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C533 N$1992 N$2361 N$1937 N$1939 "Waveguide Crossing" sch_x=58 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C534 N$2309 N$1994 N$1941 N$1943 "Waveguide Crossing" sch_x=56 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C535 N$1996 N$1998 N$1945 N$1947 "Waveguide Crossing" sch_x=56 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C536 N$2000 N$2002 N$1949 N$1951 "Waveguide Crossing" sch_x=56 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C537 N$2004 N$2006 N$1953 N$1955 "Waveguide Crossing" sch_x=56 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C538 N$2008 N$2010 N$1957 N$1959 "Waveguide Crossing" sch_x=56 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C539 N$2012 N$2014 N$1961 N$1963 "Waveguide Crossing" sch_x=56 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C540 N$2016 N$2018 N$1965 N$1967 "Waveguide Crossing" sch_x=56 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C541 N$2020 N$2022 N$1969 N$1971 "Waveguide Crossing" sch_x=56 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C542 N$2024 N$2026 N$1973 N$1975 "Waveguide Crossing" sch_x=56 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C543 N$2028 N$2030 N$1977 N$1979 "Waveguide Crossing" sch_x=56 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C544 N$2032 N$2034 N$1981 N$1983 "Waveguide Crossing" sch_x=56 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C545 N$2036 N$2038 N$1985 N$1987 "Waveguide Crossing" sch_x=56 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C546 N$2040 N$2359 N$1989 N$1991 "Waveguide Crossing" sch_x=56 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C547 N$2311 N$2042 N$1993 N$1995 "Waveguide Crossing" sch_x=54 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C548 N$2044 N$2046 N$1997 N$1999 "Waveguide Crossing" sch_x=54 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C549 N$2048 N$2050 N$2001 N$2003 "Waveguide Crossing" sch_x=54 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C550 N$2052 N$2054 N$2005 N$2007 "Waveguide Crossing" sch_x=54 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C551 N$2056 N$2058 N$2009 N$2011 "Waveguide Crossing" sch_x=54 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C552 N$2060 N$2062 N$2013 N$2015 "Waveguide Crossing" sch_x=54 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C553 N$2064 N$2066 N$2017 N$2019 "Waveguide Crossing" sch_x=54 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C554 N$2068 N$2070 N$2021 N$2023 "Waveguide Crossing" sch_x=54 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C555 N$2072 N$2074 N$2025 N$2027 "Waveguide Crossing" sch_x=54 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C556 N$2076 N$2078 N$2029 N$2031 "Waveguide Crossing" sch_x=54 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C557 N$2080 N$2082 N$2033 N$2035 "Waveguide Crossing" sch_x=54 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C558 N$2084 N$2357 N$2037 N$2039 "Waveguide Crossing" sch_x=54 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C559 N$2313 N$2086 N$2041 N$2043 "Waveguide Crossing" sch_x=52 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C560 N$2088 N$2090 N$2045 N$2047 "Waveguide Crossing" sch_x=52 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C561 N$2092 N$2094 N$2049 N$2051 "Waveguide Crossing" sch_x=52 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C562 N$2096 N$2098 N$2053 N$2055 "Waveguide Crossing" sch_x=52 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C563 N$2100 N$2102 N$2057 N$2059 "Waveguide Crossing" sch_x=52 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C564 N$2104 N$2106 N$2061 N$2063 "Waveguide Crossing" sch_x=52 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C565 N$2108 N$2110 N$2065 N$2067 "Waveguide Crossing" sch_x=52 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C566 N$2112 N$2114 N$2069 N$2071 "Waveguide Crossing" sch_x=52 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C567 N$2116 N$2118 N$2073 N$2075 "Waveguide Crossing" sch_x=52 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C568 N$2120 N$2122 N$2077 N$2079 "Waveguide Crossing" sch_x=52 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C569 N$2124 N$2355 N$2081 N$2083 "Waveguide Crossing" sch_x=52 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C570 N$2315 N$2126 N$2085 N$2087 "Waveguide Crossing" sch_x=50 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C571 N$2128 N$2130 N$2089 N$2091 "Waveguide Crossing" sch_x=50 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C572 N$2132 N$2134 N$2093 N$2095 "Waveguide Crossing" sch_x=50 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C573 N$2136 N$2138 N$2097 N$2099 "Waveguide Crossing" sch_x=50 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C574 N$2140 N$2142 N$2101 N$2103 "Waveguide Crossing" sch_x=50 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C575 N$2144 N$2146 N$2105 N$2107 "Waveguide Crossing" sch_x=50 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C576 N$2148 N$2150 N$2109 N$2111 "Waveguide Crossing" sch_x=50 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C577 N$2152 N$2154 N$2113 N$2115 "Waveguide Crossing" sch_x=50 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C578 N$2156 N$2158 N$2117 N$2119 "Waveguide Crossing" sch_x=50 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C579 N$2160 N$2353 N$2121 N$2123 "Waveguide Crossing" sch_x=50 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C580 N$2317 N$2162 N$2125 N$2127 "Waveguide Crossing" sch_x=48 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C581 N$2164 N$2166 N$2129 N$2131 "Waveguide Crossing" sch_x=48 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C582 N$2168 N$2170 N$2133 N$2135 "Waveguide Crossing" sch_x=48 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C583 N$2172 N$2174 N$2137 N$2139 "Waveguide Crossing" sch_x=48 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C584 N$2176 N$2178 N$2141 N$2143 "Waveguide Crossing" sch_x=48 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C585 N$2180 N$2182 N$2145 N$2147 "Waveguide Crossing" sch_x=48 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C586 N$2184 N$2186 N$2149 N$2151 "Waveguide Crossing" sch_x=48 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C587 N$2188 N$2190 N$2153 N$2155 "Waveguide Crossing" sch_x=48 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C588 N$2192 N$2351 N$2157 N$2159 "Waveguide Crossing" sch_x=48 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C589 N$2319 N$2194 N$2161 N$2163 "Waveguide Crossing" sch_x=46 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C590 N$2196 N$2198 N$2165 N$2167 "Waveguide Crossing" sch_x=46 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C591 N$2200 N$2202 N$2169 N$2171 "Waveguide Crossing" sch_x=46 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C592 N$2204 N$2206 N$2173 N$2175 "Waveguide Crossing" sch_x=46 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C593 N$2208 N$2210 N$2177 N$2179 "Waveguide Crossing" sch_x=46 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C594 N$2212 N$2214 N$2181 N$2183 "Waveguide Crossing" sch_x=46 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C595 N$2216 N$2218 N$2185 N$2187 "Waveguide Crossing" sch_x=46 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C596 N$2220 N$2349 N$2189 N$2191 "Waveguide Crossing" sch_x=46 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C597 N$2321 N$2222 N$2193 N$2195 "Waveguide Crossing" sch_x=44 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C598 N$2224 N$2226 N$2197 N$2199 "Waveguide Crossing" sch_x=44 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C599 N$2228 N$2230 N$2201 N$2203 "Waveguide Crossing" sch_x=44 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C600 N$2232 N$2234 N$2205 N$2207 "Waveguide Crossing" sch_x=44 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C601 N$2236 N$2238 N$2209 N$2211 "Waveguide Crossing" sch_x=44 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C602 N$2240 N$2242 N$2213 N$2215 "Waveguide Crossing" sch_x=44 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C603 N$2244 N$2347 N$2217 N$2219 "Waveguide Crossing" sch_x=44 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C604 N$2323 N$2246 N$2221 N$2223 "Waveguide Crossing" sch_x=42 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C605 N$2248 N$2250 N$2225 N$2227 "Waveguide Crossing" sch_x=42 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C606 N$2252 N$2254 N$2229 N$2231 "Waveguide Crossing" sch_x=42 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C607 N$2256 N$2258 N$2233 N$2235 "Waveguide Crossing" sch_x=42 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C608 N$2260 N$2262 N$2237 N$2239 "Waveguide Crossing" sch_x=42 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C609 N$2264 N$2345 N$2241 N$2243 "Waveguide Crossing" sch_x=42 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C610 N$2325 N$2266 N$2245 N$2247 "Waveguide Crossing" sch_x=40 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C611 N$2268 N$2270 N$2249 N$2251 "Waveguide Crossing" sch_x=40 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C612 N$2272 N$2274 N$2253 N$2255 "Waveguide Crossing" sch_x=40 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C613 N$2276 N$2278 N$2257 N$2259 "Waveguide Crossing" sch_x=40 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C614 N$2280 N$2343 N$2261 N$2263 "Waveguide Crossing" sch_x=40 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C615 N$2327 N$2282 N$2265 N$2267 "Waveguide Crossing" sch_x=38 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C616 N$2284 N$2286 N$2269 N$2271 "Waveguide Crossing" sch_x=38 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C617 N$2288 N$2290 N$2273 N$2275 "Waveguide Crossing" sch_x=38 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C618 N$2292 N$2341 N$2277 N$2279 "Waveguide Crossing" sch_x=38 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C619 N$2329 N$2294 N$2281 N$2283 "Waveguide Crossing" sch_x=36 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C620 N$2296 N$2298 N$2285 N$2287 "Waveguide Crossing" sch_x=36 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C621 N$2300 N$2339 N$2289 N$2291 "Waveguide Crossing" sch_x=36 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C622 N$2331 N$2302 N$2293 N$2295 "Waveguide Crossing" sch_x=34 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C623 N$2304 N$2337 N$2297 N$2299 "Waveguide Crossing" sch_x=34 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C624 N$2333 N$2335 N$2301 N$2303 "Waveguide Crossing" sch_x=32 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S489 N$2365 N$1826 N$8958 N$8834 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S490 N$1828 N$1830 N$8836 N$8838 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S491 N$1832 N$1834 N$8840 N$8842 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S492 N$1836 N$1838 N$8844 N$8846 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S493 N$1840 N$1842 N$8848 N$8850 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S494 N$1844 N$1846 N$8852 N$8854 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S495 N$1848 N$1850 N$8856 N$8858 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S496 N$1852 N$1854 N$8860 N$8862 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S497 N$1856 N$1858 N$8864 N$8866 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S498 N$1860 N$1862 N$8868 N$8870 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S499 N$1864 N$1866 N$8872 N$8874 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S500 N$1868 N$1870 N$8876 N$8878 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S501 N$1872 N$1874 N$8880 N$8882 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S502 N$1876 N$1878 N$8884 N$8886 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S503 N$1880 N$1882 N$8888 N$8890 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S504 N$1884 N$2367 N$8892 N$8894 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S625 N$2502 N$2490 N$2369 N$2371 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S626 N$2492 N$2494 N$2373 N$2379 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S627 N$9089 N$2370 N$2381 N$2383 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S628 N$2376 N$9090 N$2385 N$2391 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S629 N$9091 N$2378 N$2393 N$2395 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S630 N$2380 N$9092 N$2397 N$2403 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S631 N$2382 N$2390 N$2405 N$9093 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S632 N$2388 N$2392 N$9094 N$2407 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S633 N$2394 N$2402 N$2409 N$9095 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S634 N$2400 N$2404 N$9096 N$2415 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S635 N$2406 N$2414 N$2542 N$2530 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S636 N$2412 N$2416 N$2532 N$2534 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C637 N$2372 N$2374 N$2375 N$2377 "Waveguide Crossing" sch_x=-4 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C638 N$2384 N$2386 N$2389 N$2387 "Waveguide Crossing" sch_x=0 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C639 N$2396 N$2398 N$2401 N$2399 "Waveguide Crossing" sch_x=0 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C640 N$2408 N$2410 N$2413 N$2411 "Waveguide Crossing" sch_x=4 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S641 N$2496 N$2498 N$2417 N$2419 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S642 N$2500 N$2504 N$2421 N$2427 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S643 N$9097 N$2418 N$2429 N$2431 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S644 N$2424 N$9098 N$2433 N$2439 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S645 N$9099 N$2426 N$2441 N$2443 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S646 N$2428 N$9100 N$2445 N$2451 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S647 N$2430 N$2438 N$2453 N$9101 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S648 N$2436 N$2440 N$9102 N$2455 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S649 N$2442 N$2450 N$2457 N$9103 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S650 N$2448 N$2452 N$9104 N$2463 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S651 N$2454 N$2462 N$2536 N$2538 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S652 N$2460 N$2464 N$2540 N$2544 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C653 N$2420 N$2422 N$2423 N$2425 "Waveguide Crossing" sch_x=-4 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C654 N$2432 N$2434 N$2437 N$2435 "Waveguide Crossing" sch_x=0 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C655 N$2444 N$2446 N$2449 N$2447 "Waveguide Crossing" sch_x=0 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C656 N$2456 N$2458 N$2461 N$2459 "Waveguide Crossing" sch_x=4 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C671 N$2529 N$2518 N$2505 N$2507 "Waveguide Crossing" sch_x=12 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C672 N$2520 N$2522 N$2509 N$2511 "Waveguide Crossing" sch_x=12 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C673 N$2524 N$2539 N$2513 N$2515 "Waveguide Crossing" sch_x=12 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C674 N$2531 N$2526 N$2517 N$2519 "Waveguide Crossing" sch_x=10 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C675 N$2528 N$2537 N$2521 N$2523 "Waveguide Crossing" sch_x=10 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C676 N$2533 N$2535 N$2525 N$2527 "Waveguide Crossing" sch_x=8 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S667 N$2541 N$2506 N$3006 N$2978 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S668 N$2508 N$2510 N$2980 N$2982 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S669 N$2512 N$2514 N$2984 N$2986 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S670 N$2516 N$2543 N$2988 N$2990 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S677 N$2678 N$2666 N$2545 N$2547 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S678 N$2668 N$2670 N$2549 N$2555 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S679 N$9105 N$2546 N$2557 N$2559 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S680 N$2552 N$9106 N$2561 N$2567 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S681 N$9107 N$2554 N$2569 N$2571 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S682 N$2556 N$9108 N$2573 N$2579 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S683 N$2558 N$2566 N$2581 N$9109 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S684 N$2564 N$2568 N$9110 N$2583 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S685 N$2570 N$2578 N$2585 N$9111 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S686 N$2576 N$2580 N$9112 N$2591 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S687 N$2582 N$2590 N$2718 N$2706 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S688 N$2588 N$2592 N$2708 N$2710 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C689 N$2548 N$2550 N$2551 N$2553 "Waveguide Crossing" sch_x=-4 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C690 N$2560 N$2562 N$2565 N$2563 "Waveguide Crossing" sch_x=0 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C691 N$2572 N$2574 N$2577 N$2575 "Waveguide Crossing" sch_x=0 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C692 N$2584 N$2586 N$2589 N$2587 "Waveguide Crossing" sch_x=4 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S693 N$2672 N$2674 N$2593 N$2595 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S694 N$2676 N$2680 N$2597 N$2603 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S695 N$9113 N$2594 N$2605 N$2607 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S696 N$2600 N$9114 N$2609 N$2615 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S697 N$9115 N$2602 N$2617 N$2619 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S698 N$2604 N$9116 N$2621 N$2627 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S699 N$2606 N$2614 N$2629 N$9117 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S700 N$2612 N$2616 N$9118 N$2631 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S701 N$2618 N$2626 N$2633 N$9119 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S702 N$2624 N$2628 N$9120 N$2639 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S703 N$2630 N$2638 N$2712 N$2714 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S704 N$2636 N$2640 N$2716 N$2720 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C705 N$2596 N$2598 N$2599 N$2601 "Waveguide Crossing" sch_x=-4 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C706 N$2608 N$2610 N$2613 N$2611 "Waveguide Crossing" sch_x=0 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C707 N$2620 N$2622 N$2625 N$2623 "Waveguide Crossing" sch_x=0 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C708 N$2632 N$2634 N$2637 N$2635 "Waveguide Crossing" sch_x=4 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C723 N$2705 N$2694 N$2681 N$2683 "Waveguide Crossing" sch_x=12 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C724 N$2696 N$2698 N$2685 N$2687 "Waveguide Crossing" sch_x=12 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C725 N$2700 N$2715 N$2689 N$2691 "Waveguide Crossing" sch_x=12 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C726 N$2707 N$2702 N$2693 N$2695 "Waveguide Crossing" sch_x=10 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C727 N$2704 N$2713 N$2697 N$2699 "Waveguide Crossing" sch_x=10 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C728 N$2709 N$2711 N$2701 N$2703 "Waveguide Crossing" sch_x=8 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S719 N$2717 N$2682 N$2992 N$2994 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S720 N$2684 N$2686 N$2996 N$2998 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S721 N$2688 N$2690 N$3000 N$3002 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S722 N$2692 N$2719 N$3004 N$3008 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C773 N$2977 N$2894 N$2865 N$2867 "Waveguide Crossing" sch_x=28 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C774 N$2896 N$2898 N$2869 N$2871 "Waveguide Crossing" sch_x=28 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C775 N$2900 N$2902 N$2873 N$2875 "Waveguide Crossing" sch_x=28 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C776 N$2904 N$2906 N$2877 N$2879 "Waveguide Crossing" sch_x=28 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C777 N$2908 N$2910 N$2881 N$2883 "Waveguide Crossing" sch_x=28 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C778 N$2912 N$2914 N$2885 N$2887 "Waveguide Crossing" sch_x=28 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C779 N$2916 N$3003 N$2889 N$2891 "Waveguide Crossing" sch_x=28 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C780 N$2979 N$2918 N$2893 N$2895 "Waveguide Crossing" sch_x=26 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C781 N$2920 N$2922 N$2897 N$2899 "Waveguide Crossing" sch_x=26 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C782 N$2924 N$2926 N$2901 N$2903 "Waveguide Crossing" sch_x=26 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C783 N$2928 N$2930 N$2905 N$2907 "Waveguide Crossing" sch_x=26 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C784 N$2932 N$2934 N$2909 N$2911 "Waveguide Crossing" sch_x=26 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C785 N$2936 N$3001 N$2913 N$2915 "Waveguide Crossing" sch_x=26 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C786 N$2981 N$2938 N$2917 N$2919 "Waveguide Crossing" sch_x=24 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C787 N$2940 N$2942 N$2921 N$2923 "Waveguide Crossing" sch_x=24 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C788 N$2944 N$2946 N$2925 N$2927 "Waveguide Crossing" sch_x=24 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C789 N$2948 N$2950 N$2929 N$2931 "Waveguide Crossing" sch_x=24 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C790 N$2952 N$2999 N$2933 N$2935 "Waveguide Crossing" sch_x=24 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C791 N$2983 N$2954 N$2937 N$2939 "Waveguide Crossing" sch_x=22 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C792 N$2956 N$2958 N$2941 N$2943 "Waveguide Crossing" sch_x=22 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C793 N$2960 N$2962 N$2945 N$2947 "Waveguide Crossing" sch_x=22 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C794 N$2964 N$2997 N$2949 N$2951 "Waveguide Crossing" sch_x=22 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C795 N$2985 N$2966 N$2953 N$2955 "Waveguide Crossing" sch_x=20 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C796 N$2968 N$2970 N$2957 N$2959 "Waveguide Crossing" sch_x=20 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C797 N$2972 N$2995 N$2961 N$2963 "Waveguide Crossing" sch_x=20 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C798 N$2987 N$2974 N$2965 N$2967 "Waveguide Crossing" sch_x=18 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C799 N$2976 N$2993 N$2969 N$2971 "Waveguide Crossing" sch_x=18 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C800 N$2989 N$2991 N$2973 N$2975 "Waveguide Crossing" sch_x=16 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S765 N$3005 N$2866 N$4734 N$4674 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S766 N$2868 N$2870 N$4676 N$4678 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S767 N$2872 N$2874 N$4680 N$4682 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S768 N$2876 N$2878 N$4684 N$4686 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S769 N$2880 N$2882 N$4688 N$4690 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S770 N$2884 N$2886 N$4692 N$4694 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S771 N$2888 N$2890 N$4696 N$4698 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S772 N$2892 N$3007 N$4700 N$4702 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S801 N$3142 N$3130 N$3009 N$3011 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S802 N$3132 N$3134 N$3013 N$3019 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S803 N$9121 N$3010 N$3021 N$3023 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S804 N$3016 N$9122 N$3025 N$3031 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S805 N$9123 N$3018 N$3033 N$3035 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S806 N$3020 N$9124 N$3037 N$3043 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S807 N$3022 N$3030 N$3045 N$9125 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S808 N$3028 N$3032 N$9126 N$3047 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S809 N$3034 N$3042 N$3049 N$9127 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S810 N$3040 N$3044 N$9128 N$3055 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S811 N$3046 N$3054 N$3182 N$3170 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S812 N$3052 N$3056 N$3172 N$3174 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C813 N$3012 N$3014 N$3015 N$3017 "Waveguide Crossing" sch_x=-4 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C814 N$3024 N$3026 N$3029 N$3027 "Waveguide Crossing" sch_x=0 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C815 N$3036 N$3038 N$3041 N$3039 "Waveguide Crossing" sch_x=0 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C816 N$3048 N$3050 N$3053 N$3051 "Waveguide Crossing" sch_x=4 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S817 N$3136 N$3138 N$3057 N$3059 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S818 N$3140 N$3144 N$3061 N$3067 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S819 N$9129 N$3058 N$3069 N$3071 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S820 N$3064 N$9130 N$3073 N$3079 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S821 N$9131 N$3066 N$3081 N$3083 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S822 N$3068 N$9132 N$3085 N$3091 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S823 N$3070 N$3078 N$3093 N$9133 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S824 N$3076 N$3080 N$9134 N$3095 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S825 N$3082 N$3090 N$3097 N$9135 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S826 N$3088 N$3092 N$9136 N$3103 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S827 N$3094 N$3102 N$3176 N$3178 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S828 N$3100 N$3104 N$3180 N$3184 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C829 N$3060 N$3062 N$3063 N$3065 "Waveguide Crossing" sch_x=-4 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C830 N$3072 N$3074 N$3077 N$3075 "Waveguide Crossing" sch_x=0 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C831 N$3084 N$3086 N$3089 N$3087 "Waveguide Crossing" sch_x=0 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C832 N$3096 N$3098 N$3101 N$3099 "Waveguide Crossing" sch_x=4 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C847 N$3169 N$3158 N$3145 N$3147 "Waveguide Crossing" sch_x=12 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C848 N$3160 N$3162 N$3149 N$3151 "Waveguide Crossing" sch_x=12 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C849 N$3164 N$3179 N$3153 N$3155 "Waveguide Crossing" sch_x=12 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C850 N$3171 N$3166 N$3157 N$3159 "Waveguide Crossing" sch_x=10 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C851 N$3168 N$3177 N$3161 N$3163 "Waveguide Crossing" sch_x=10 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C852 N$3173 N$3175 N$3165 N$3167 "Waveguide Crossing" sch_x=8 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S843 N$3181 N$3146 N$3646 N$3618 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S844 N$3148 N$3150 N$3620 N$3622 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S845 N$3152 N$3154 N$3624 N$3626 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S846 N$3156 N$3183 N$3628 N$3630 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S853 N$3318 N$3306 N$3185 N$3187 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S854 N$3308 N$3310 N$3189 N$3195 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S855 N$9137 N$3186 N$3197 N$3199 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S856 N$3192 N$9138 N$3201 N$3207 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S857 N$9139 N$3194 N$3209 N$3211 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S858 N$3196 N$9140 N$3213 N$3219 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S859 N$3198 N$3206 N$3221 N$9141 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S860 N$3204 N$3208 N$9142 N$3223 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S861 N$3210 N$3218 N$3225 N$9143 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S862 N$3216 N$3220 N$9144 N$3231 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S863 N$3222 N$3230 N$3358 N$3346 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S864 N$3228 N$3232 N$3348 N$3350 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C865 N$3188 N$3190 N$3191 N$3193 "Waveguide Crossing" sch_x=-4 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C866 N$3200 N$3202 N$3205 N$3203 "Waveguide Crossing" sch_x=0 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C867 N$3212 N$3214 N$3217 N$3215 "Waveguide Crossing" sch_x=0 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C868 N$3224 N$3226 N$3229 N$3227 "Waveguide Crossing" sch_x=4 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S869 N$3312 N$3314 N$3233 N$3235 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S870 N$3316 N$3320 N$3237 N$3243 MMI_switch_ideal library="Design kits/capstone" sch_x=-6 sch_y=-30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S871 N$9145 N$3234 N$3245 N$3247 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S872 N$3240 N$9146 N$3249 N$3255 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S873 N$9147 N$3242 N$3257 N$3259 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S874 N$3244 N$9148 N$3261 N$3267 MMI_switch_ideal library="Design kits/capstone" sch_x=-2 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S875 N$3246 N$3254 N$3269 N$9149 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S876 N$3252 N$3256 N$9150 N$3271 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S877 N$3258 N$3266 N$3273 N$9151 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S878 N$3264 N$3268 N$9152 N$3279 MMI_switch_ideal library="Design kits/capstone" sch_x=2 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S879 N$3270 N$3278 N$3352 N$3354 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S880 N$3276 N$3280 N$3356 N$3360 MMI_switch_ideal library="Design kits/capstone" sch_x=6 sch_y=-30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C881 N$3236 N$3238 N$3239 N$3241 "Waveguide Crossing" sch_x=-4 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C882 N$3248 N$3250 N$3253 N$3251 "Waveguide Crossing" sch_x=0 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C883 N$3260 N$3262 N$3265 N$3263 "Waveguide Crossing" sch_x=0 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C884 N$3272 N$3274 N$3277 N$3275 "Waveguide Crossing" sch_x=4 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C899 N$3345 N$3334 N$3321 N$3323 "Waveguide Crossing" sch_x=12 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C900 N$3336 N$3338 N$3325 N$3327 "Waveguide Crossing" sch_x=12 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C901 N$3340 N$3355 N$3329 N$3331 "Waveguide Crossing" sch_x=12 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C902 N$3347 N$3342 N$3333 N$3335 "Waveguide Crossing" sch_x=10 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C903 N$3344 N$3353 N$3337 N$3339 "Waveguide Crossing" sch_x=10 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C904 N$3349 N$3351 N$3341 N$3343 "Waveguide Crossing" sch_x=8 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S895 N$3357 N$3322 N$3632 N$3634 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S896 N$3324 N$3326 N$3636 N$3638 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S897 N$3328 N$3330 N$3640 N$3642 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S898 N$3332 N$3359 N$3644 N$3648 MMI_switch_ideal library="Design kits/capstone" sch_x=14 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C949 N$3617 N$3534 N$3505 N$3507 "Waveguide Crossing" sch_x=28 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C950 N$3536 N$3538 N$3509 N$3511 "Waveguide Crossing" sch_x=28 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C951 N$3540 N$3542 N$3513 N$3515 "Waveguide Crossing" sch_x=28 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C952 N$3544 N$3546 N$3517 N$3519 "Waveguide Crossing" sch_x=28 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C953 N$3548 N$3550 N$3521 N$3523 "Waveguide Crossing" sch_x=28 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C954 N$3552 N$3554 N$3525 N$3527 "Waveguide Crossing" sch_x=28 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C955 N$3556 N$3643 N$3529 N$3531 "Waveguide Crossing" sch_x=28 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C956 N$3619 N$3558 N$3533 N$3535 "Waveguide Crossing" sch_x=26 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C957 N$3560 N$3562 N$3537 N$3539 "Waveguide Crossing" sch_x=26 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C958 N$3564 N$3566 N$3541 N$3543 "Waveguide Crossing" sch_x=26 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C959 N$3568 N$3570 N$3545 N$3547 "Waveguide Crossing" sch_x=26 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C960 N$3572 N$3574 N$3549 N$3551 "Waveguide Crossing" sch_x=26 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C961 N$3576 N$3641 N$3553 N$3555 "Waveguide Crossing" sch_x=26 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C962 N$3621 N$3578 N$3557 N$3559 "Waveguide Crossing" sch_x=24 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C963 N$3580 N$3582 N$3561 N$3563 "Waveguide Crossing" sch_x=24 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C964 N$3584 N$3586 N$3565 N$3567 "Waveguide Crossing" sch_x=24 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C965 N$3588 N$3590 N$3569 N$3571 "Waveguide Crossing" sch_x=24 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C966 N$3592 N$3639 N$3573 N$3575 "Waveguide Crossing" sch_x=24 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C967 N$3623 N$3594 N$3577 N$3579 "Waveguide Crossing" sch_x=22 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C968 N$3596 N$3598 N$3581 N$3583 "Waveguide Crossing" sch_x=22 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C969 N$3600 N$3602 N$3585 N$3587 "Waveguide Crossing" sch_x=22 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C970 N$3604 N$3637 N$3589 N$3591 "Waveguide Crossing" sch_x=22 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C971 N$3625 N$3606 N$3593 N$3595 "Waveguide Crossing" sch_x=20 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C972 N$3608 N$3610 N$3597 N$3599 "Waveguide Crossing" sch_x=20 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C973 N$3612 N$3635 N$3601 N$3603 "Waveguide Crossing" sch_x=20 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C974 N$3627 N$3614 N$3605 N$3607 "Waveguide Crossing" sch_x=18 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C975 N$3616 N$3633 N$3609 N$3611 "Waveguide Crossing" sch_x=18 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C976 N$3629 N$3631 N$3613 N$3615 "Waveguide Crossing" sch_x=16 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S941 N$3645 N$3506 N$4704 N$4706 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S942 N$3508 N$3510 N$4708 N$4710 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S943 N$3512 N$3514 N$4712 N$4714 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S944 N$3516 N$3518 N$4716 N$4718 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S945 N$3520 N$3522 N$4720 N$4722 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S946 N$3524 N$3526 N$4724 N$4726 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S947 N$3528 N$3530 N$4728 N$4730 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S948 N$3532 N$3647 N$4732 N$4736 MMI_switch_ideal library="Design kits/capstone" sch_x=30 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1129 N$4673 N$4254 N$4193 N$4195 "Waveguide Crossing" sch_x=60 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1130 N$4256 N$4258 N$4197 N$4199 "Waveguide Crossing" sch_x=60 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1131 N$4260 N$4262 N$4201 N$4203 "Waveguide Crossing" sch_x=60 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1132 N$4264 N$4266 N$4205 N$4207 "Waveguide Crossing" sch_x=60 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1133 N$4268 N$4270 N$4209 N$4211 "Waveguide Crossing" sch_x=60 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1134 N$4272 N$4274 N$4213 N$4215 "Waveguide Crossing" sch_x=60 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1135 N$4276 N$4278 N$4217 N$4219 "Waveguide Crossing" sch_x=60 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1136 N$4280 N$4282 N$4221 N$4223 "Waveguide Crossing" sch_x=60 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1137 N$4284 N$4286 N$4225 N$4227 "Waveguide Crossing" sch_x=60 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1138 N$4288 N$4290 N$4229 N$4231 "Waveguide Crossing" sch_x=60 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1139 N$4292 N$4294 N$4233 N$4235 "Waveguide Crossing" sch_x=60 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1140 N$4296 N$4298 N$4237 N$4239 "Waveguide Crossing" sch_x=60 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1141 N$4300 N$4302 N$4241 N$4243 "Waveguide Crossing" sch_x=60 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1142 N$4304 N$4306 N$4245 N$4247 "Waveguide Crossing" sch_x=60 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1143 N$4308 N$4731 N$4249 N$4251 "Waveguide Crossing" sch_x=60 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1144 N$4675 N$4310 N$4253 N$4255 "Waveguide Crossing" sch_x=58 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1145 N$4312 N$4314 N$4257 N$4259 "Waveguide Crossing" sch_x=58 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1146 N$4316 N$4318 N$4261 N$4263 "Waveguide Crossing" sch_x=58 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1147 N$4320 N$4322 N$4265 N$4267 "Waveguide Crossing" sch_x=58 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1148 N$4324 N$4326 N$4269 N$4271 "Waveguide Crossing" sch_x=58 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1149 N$4328 N$4330 N$4273 N$4275 "Waveguide Crossing" sch_x=58 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1150 N$4332 N$4334 N$4277 N$4279 "Waveguide Crossing" sch_x=58 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1151 N$4336 N$4338 N$4281 N$4283 "Waveguide Crossing" sch_x=58 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1152 N$4340 N$4342 N$4285 N$4287 "Waveguide Crossing" sch_x=58 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1153 N$4344 N$4346 N$4289 N$4291 "Waveguide Crossing" sch_x=58 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1154 N$4348 N$4350 N$4293 N$4295 "Waveguide Crossing" sch_x=58 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1155 N$4352 N$4354 N$4297 N$4299 "Waveguide Crossing" sch_x=58 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1156 N$4356 N$4358 N$4301 N$4303 "Waveguide Crossing" sch_x=58 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1157 N$4360 N$4729 N$4305 N$4307 "Waveguide Crossing" sch_x=58 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1158 N$4677 N$4362 N$4309 N$4311 "Waveguide Crossing" sch_x=56 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1159 N$4364 N$4366 N$4313 N$4315 "Waveguide Crossing" sch_x=56 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1160 N$4368 N$4370 N$4317 N$4319 "Waveguide Crossing" sch_x=56 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1161 N$4372 N$4374 N$4321 N$4323 "Waveguide Crossing" sch_x=56 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1162 N$4376 N$4378 N$4325 N$4327 "Waveguide Crossing" sch_x=56 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1163 N$4380 N$4382 N$4329 N$4331 "Waveguide Crossing" sch_x=56 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1164 N$4384 N$4386 N$4333 N$4335 "Waveguide Crossing" sch_x=56 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1165 N$4388 N$4390 N$4337 N$4339 "Waveguide Crossing" sch_x=56 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1166 N$4392 N$4394 N$4341 N$4343 "Waveguide Crossing" sch_x=56 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1167 N$4396 N$4398 N$4345 N$4347 "Waveguide Crossing" sch_x=56 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1168 N$4400 N$4402 N$4349 N$4351 "Waveguide Crossing" sch_x=56 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1169 N$4404 N$4406 N$4353 N$4355 "Waveguide Crossing" sch_x=56 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1170 N$4408 N$4727 N$4357 N$4359 "Waveguide Crossing" sch_x=56 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1171 N$4679 N$4410 N$4361 N$4363 "Waveguide Crossing" sch_x=54 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1172 N$4412 N$4414 N$4365 N$4367 "Waveguide Crossing" sch_x=54 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1173 N$4416 N$4418 N$4369 N$4371 "Waveguide Crossing" sch_x=54 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1174 N$4420 N$4422 N$4373 N$4375 "Waveguide Crossing" sch_x=54 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1175 N$4424 N$4426 N$4377 N$4379 "Waveguide Crossing" sch_x=54 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1176 N$4428 N$4430 N$4381 N$4383 "Waveguide Crossing" sch_x=54 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1177 N$4432 N$4434 N$4385 N$4387 "Waveguide Crossing" sch_x=54 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1178 N$4436 N$4438 N$4389 N$4391 "Waveguide Crossing" sch_x=54 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1179 N$4440 N$4442 N$4393 N$4395 "Waveguide Crossing" sch_x=54 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1180 N$4444 N$4446 N$4397 N$4399 "Waveguide Crossing" sch_x=54 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1181 N$4448 N$4450 N$4401 N$4403 "Waveguide Crossing" sch_x=54 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1182 N$4452 N$4725 N$4405 N$4407 "Waveguide Crossing" sch_x=54 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1183 N$4681 N$4454 N$4409 N$4411 "Waveguide Crossing" sch_x=52 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1184 N$4456 N$4458 N$4413 N$4415 "Waveguide Crossing" sch_x=52 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1185 N$4460 N$4462 N$4417 N$4419 "Waveguide Crossing" sch_x=52 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1186 N$4464 N$4466 N$4421 N$4423 "Waveguide Crossing" sch_x=52 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1187 N$4468 N$4470 N$4425 N$4427 "Waveguide Crossing" sch_x=52 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1188 N$4472 N$4474 N$4429 N$4431 "Waveguide Crossing" sch_x=52 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1189 N$4476 N$4478 N$4433 N$4435 "Waveguide Crossing" sch_x=52 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1190 N$4480 N$4482 N$4437 N$4439 "Waveguide Crossing" sch_x=52 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1191 N$4484 N$4486 N$4441 N$4443 "Waveguide Crossing" sch_x=52 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1192 N$4488 N$4490 N$4445 N$4447 "Waveguide Crossing" sch_x=52 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1193 N$4492 N$4723 N$4449 N$4451 "Waveguide Crossing" sch_x=52 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1194 N$4683 N$4494 N$4453 N$4455 "Waveguide Crossing" sch_x=50 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1195 N$4496 N$4498 N$4457 N$4459 "Waveguide Crossing" sch_x=50 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1196 N$4500 N$4502 N$4461 N$4463 "Waveguide Crossing" sch_x=50 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1197 N$4504 N$4506 N$4465 N$4467 "Waveguide Crossing" sch_x=50 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1198 N$4508 N$4510 N$4469 N$4471 "Waveguide Crossing" sch_x=50 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1199 N$4512 N$4514 N$4473 N$4475 "Waveguide Crossing" sch_x=50 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1200 N$4516 N$4518 N$4477 N$4479 "Waveguide Crossing" sch_x=50 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1201 N$4520 N$4522 N$4481 N$4483 "Waveguide Crossing" sch_x=50 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1202 N$4524 N$4526 N$4485 N$4487 "Waveguide Crossing" sch_x=50 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1203 N$4528 N$4721 N$4489 N$4491 "Waveguide Crossing" sch_x=50 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1204 N$4685 N$4530 N$4493 N$4495 "Waveguide Crossing" sch_x=48 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1205 N$4532 N$4534 N$4497 N$4499 "Waveguide Crossing" sch_x=48 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1206 N$4536 N$4538 N$4501 N$4503 "Waveguide Crossing" sch_x=48 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1207 N$4540 N$4542 N$4505 N$4507 "Waveguide Crossing" sch_x=48 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1208 N$4544 N$4546 N$4509 N$4511 "Waveguide Crossing" sch_x=48 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1209 N$4548 N$4550 N$4513 N$4515 "Waveguide Crossing" sch_x=48 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1210 N$4552 N$4554 N$4517 N$4519 "Waveguide Crossing" sch_x=48 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1211 N$4556 N$4558 N$4521 N$4523 "Waveguide Crossing" sch_x=48 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1212 N$4560 N$4719 N$4525 N$4527 "Waveguide Crossing" sch_x=48 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1213 N$4687 N$4562 N$4529 N$4531 "Waveguide Crossing" sch_x=46 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1214 N$4564 N$4566 N$4533 N$4535 "Waveguide Crossing" sch_x=46 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1215 N$4568 N$4570 N$4537 N$4539 "Waveguide Crossing" sch_x=46 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1216 N$4572 N$4574 N$4541 N$4543 "Waveguide Crossing" sch_x=46 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1217 N$4576 N$4578 N$4545 N$4547 "Waveguide Crossing" sch_x=46 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1218 N$4580 N$4582 N$4549 N$4551 "Waveguide Crossing" sch_x=46 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1219 N$4584 N$4586 N$4553 N$4555 "Waveguide Crossing" sch_x=46 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1220 N$4588 N$4717 N$4557 N$4559 "Waveguide Crossing" sch_x=46 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1221 N$4689 N$4590 N$4561 N$4563 "Waveguide Crossing" sch_x=44 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1222 N$4592 N$4594 N$4565 N$4567 "Waveguide Crossing" sch_x=44 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1223 N$4596 N$4598 N$4569 N$4571 "Waveguide Crossing" sch_x=44 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1224 N$4600 N$4602 N$4573 N$4575 "Waveguide Crossing" sch_x=44 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1225 N$4604 N$4606 N$4577 N$4579 "Waveguide Crossing" sch_x=44 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1226 N$4608 N$4610 N$4581 N$4583 "Waveguide Crossing" sch_x=44 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1227 N$4612 N$4715 N$4585 N$4587 "Waveguide Crossing" sch_x=44 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1228 N$4691 N$4614 N$4589 N$4591 "Waveguide Crossing" sch_x=42 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1229 N$4616 N$4618 N$4593 N$4595 "Waveguide Crossing" sch_x=42 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1230 N$4620 N$4622 N$4597 N$4599 "Waveguide Crossing" sch_x=42 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1231 N$4624 N$4626 N$4601 N$4603 "Waveguide Crossing" sch_x=42 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1232 N$4628 N$4630 N$4605 N$4607 "Waveguide Crossing" sch_x=42 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1233 N$4632 N$4713 N$4609 N$4611 "Waveguide Crossing" sch_x=42 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1234 N$4693 N$4634 N$4613 N$4615 "Waveguide Crossing" sch_x=40 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1235 N$4636 N$4638 N$4617 N$4619 "Waveguide Crossing" sch_x=40 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1236 N$4640 N$4642 N$4621 N$4623 "Waveguide Crossing" sch_x=40 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1237 N$4644 N$4646 N$4625 N$4627 "Waveguide Crossing" sch_x=40 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1238 N$4648 N$4711 N$4629 N$4631 "Waveguide Crossing" sch_x=40 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1239 N$4695 N$4650 N$4633 N$4635 "Waveguide Crossing" sch_x=38 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1240 N$4652 N$4654 N$4637 N$4639 "Waveguide Crossing" sch_x=38 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1241 N$4656 N$4658 N$4641 N$4643 "Waveguide Crossing" sch_x=38 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1242 N$4660 N$4709 N$4645 N$4647 "Waveguide Crossing" sch_x=38 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1243 N$4697 N$4662 N$4649 N$4651 "Waveguide Crossing" sch_x=36 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1244 N$4664 N$4666 N$4653 N$4655 "Waveguide Crossing" sch_x=36 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1245 N$4668 N$4707 N$4657 N$4659 "Waveguide Crossing" sch_x=36 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1246 N$4699 N$4670 N$4661 N$4663 "Waveguide Crossing" sch_x=34 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1247 N$4672 N$4705 N$4665 N$4667 "Waveguide Crossing" sch_x=34 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1248 N$4701 N$4703 N$4669 N$4671 "Waveguide Crossing" sch_x=32 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1113 N$4733 N$4194 N$8896 N$8898 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1114 N$4196 N$4198 N$8900 N$8902 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1115 N$4200 N$4202 N$8904 N$8906 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1116 N$4204 N$4206 N$8908 N$8910 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1117 N$4208 N$4210 N$8912 N$8914 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1118 N$4212 N$4214 N$8916 N$8918 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1119 N$4216 N$4218 N$8920 N$8922 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1120 N$4220 N$4222 N$8924 N$8926 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1121 N$4224 N$4226 N$8928 N$8930 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1122 N$4228 N$4230 N$8932 N$8934 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1123 N$4232 N$4234 N$8936 N$8938 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1124 N$4236 N$4238 N$8940 N$8942 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1125 N$4240 N$4242 N$8944 N$8946 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1126 N$4244 N$4246 N$8948 N$8950 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1127 N$4248 N$4250 N$8952 N$8954 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1128 N$4252 N$4735 N$8956 N$8960 MMI_switch_ideal library="Design kits/capstone" sch_x=62 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1809 N$8833 N$6974 N$6849 N$6851 "Waveguide Crossing" sch_x=124 sch_y=30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1810 N$6976 N$6978 N$6853 N$6855 "Waveguide Crossing" sch_x=124 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1811 N$6980 N$6982 N$6857 N$6859 "Waveguide Crossing" sch_x=124 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1812 N$6984 N$6986 N$6861 N$6863 "Waveguide Crossing" sch_x=124 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1813 N$6988 N$6990 N$6865 N$6867 "Waveguide Crossing" sch_x=124 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1814 N$6992 N$6994 N$6869 N$6871 "Waveguide Crossing" sch_x=124 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1815 N$6996 N$6998 N$6873 N$6875 "Waveguide Crossing" sch_x=124 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1816 N$7000 N$7002 N$6877 N$6879 "Waveguide Crossing" sch_x=124 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1817 N$7004 N$7006 N$6881 N$6883 "Waveguide Crossing" sch_x=124 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1818 N$7008 N$7010 N$6885 N$6887 "Waveguide Crossing" sch_x=124 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1819 N$7012 N$7014 N$6889 N$6891 "Waveguide Crossing" sch_x=124 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1820 N$7016 N$7018 N$6893 N$6895 "Waveguide Crossing" sch_x=124 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1821 N$7020 N$7022 N$6897 N$6899 "Waveguide Crossing" sch_x=124 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1822 N$7024 N$7026 N$6901 N$6903 "Waveguide Crossing" sch_x=124 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1823 N$7028 N$7030 N$6905 N$6907 "Waveguide Crossing" sch_x=124 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1824 N$7032 N$7034 N$6909 N$6911 "Waveguide Crossing" sch_x=124 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1825 N$7036 N$7038 N$6913 N$6915 "Waveguide Crossing" sch_x=124 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1826 N$7040 N$7042 N$6917 N$6919 "Waveguide Crossing" sch_x=124 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1827 N$7044 N$7046 N$6921 N$6923 "Waveguide Crossing" sch_x=124 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1828 N$7048 N$7050 N$6925 N$6927 "Waveguide Crossing" sch_x=124 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1829 N$7052 N$7054 N$6929 N$6931 "Waveguide Crossing" sch_x=124 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1830 N$7056 N$7058 N$6933 N$6935 "Waveguide Crossing" sch_x=124 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1831 N$7060 N$7062 N$6937 N$6939 "Waveguide Crossing" sch_x=124 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1832 N$7064 N$7066 N$6941 N$6943 "Waveguide Crossing" sch_x=124 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1833 N$7068 N$7070 N$6945 N$6947 "Waveguide Crossing" sch_x=124 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1834 N$7072 N$7074 N$6949 N$6951 "Waveguide Crossing" sch_x=124 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1835 N$7076 N$7078 N$6953 N$6955 "Waveguide Crossing" sch_x=124 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1836 N$7080 N$7082 N$6957 N$6959 "Waveguide Crossing" sch_x=124 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1837 N$7084 N$7086 N$6961 N$6963 "Waveguide Crossing" sch_x=124 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1838 N$7088 N$7090 N$6965 N$6967 "Waveguide Crossing" sch_x=124 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1839 N$7092 N$8955 N$6969 N$6971 "Waveguide Crossing" sch_x=124 sch_y=-30 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1840 N$8835 N$7094 N$6973 N$6975 "Waveguide Crossing" sch_x=122 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1841 N$7096 N$7098 N$6977 N$6979 "Waveguide Crossing" sch_x=122 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1842 N$7100 N$7102 N$6981 N$6983 "Waveguide Crossing" sch_x=122 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1843 N$7104 N$7106 N$6985 N$6987 "Waveguide Crossing" sch_x=122 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1844 N$7108 N$7110 N$6989 N$6991 "Waveguide Crossing" sch_x=122 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1845 N$7112 N$7114 N$6993 N$6995 "Waveguide Crossing" sch_x=122 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1846 N$7116 N$7118 N$6997 N$6999 "Waveguide Crossing" sch_x=122 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1847 N$7120 N$7122 N$7001 N$7003 "Waveguide Crossing" sch_x=122 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1848 N$7124 N$7126 N$7005 N$7007 "Waveguide Crossing" sch_x=122 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1849 N$7128 N$7130 N$7009 N$7011 "Waveguide Crossing" sch_x=122 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1850 N$7132 N$7134 N$7013 N$7015 "Waveguide Crossing" sch_x=122 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1851 N$7136 N$7138 N$7017 N$7019 "Waveguide Crossing" sch_x=122 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1852 N$7140 N$7142 N$7021 N$7023 "Waveguide Crossing" sch_x=122 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1853 N$7144 N$7146 N$7025 N$7027 "Waveguide Crossing" sch_x=122 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1854 N$7148 N$7150 N$7029 N$7031 "Waveguide Crossing" sch_x=122 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1855 N$7152 N$7154 N$7033 N$7035 "Waveguide Crossing" sch_x=122 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1856 N$7156 N$7158 N$7037 N$7039 "Waveguide Crossing" sch_x=122 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1857 N$7160 N$7162 N$7041 N$7043 "Waveguide Crossing" sch_x=122 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1858 N$7164 N$7166 N$7045 N$7047 "Waveguide Crossing" sch_x=122 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1859 N$7168 N$7170 N$7049 N$7051 "Waveguide Crossing" sch_x=122 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1860 N$7172 N$7174 N$7053 N$7055 "Waveguide Crossing" sch_x=122 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1861 N$7176 N$7178 N$7057 N$7059 "Waveguide Crossing" sch_x=122 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1862 N$7180 N$7182 N$7061 N$7063 "Waveguide Crossing" sch_x=122 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1863 N$7184 N$7186 N$7065 N$7067 "Waveguide Crossing" sch_x=122 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1864 N$7188 N$7190 N$7069 N$7071 "Waveguide Crossing" sch_x=122 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1865 N$7192 N$7194 N$7073 N$7075 "Waveguide Crossing" sch_x=122 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1866 N$7196 N$7198 N$7077 N$7079 "Waveguide Crossing" sch_x=122 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1867 N$7200 N$7202 N$7081 N$7083 "Waveguide Crossing" sch_x=122 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1868 N$7204 N$7206 N$7085 N$7087 "Waveguide Crossing" sch_x=122 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1869 N$7208 N$8953 N$7089 N$7091 "Waveguide Crossing" sch_x=122 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1870 N$8837 N$7210 N$7093 N$7095 "Waveguide Crossing" sch_x=120 sch_y=28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1871 N$7212 N$7214 N$7097 N$7099 "Waveguide Crossing" sch_x=120 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1872 N$7216 N$7218 N$7101 N$7103 "Waveguide Crossing" sch_x=120 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1873 N$7220 N$7222 N$7105 N$7107 "Waveguide Crossing" sch_x=120 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1874 N$7224 N$7226 N$7109 N$7111 "Waveguide Crossing" sch_x=120 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1875 N$7228 N$7230 N$7113 N$7115 "Waveguide Crossing" sch_x=120 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1876 N$7232 N$7234 N$7117 N$7119 "Waveguide Crossing" sch_x=120 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1877 N$7236 N$7238 N$7121 N$7123 "Waveguide Crossing" sch_x=120 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1878 N$7240 N$7242 N$7125 N$7127 "Waveguide Crossing" sch_x=120 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1879 N$7244 N$7246 N$7129 N$7131 "Waveguide Crossing" sch_x=120 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1880 N$7248 N$7250 N$7133 N$7135 "Waveguide Crossing" sch_x=120 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1881 N$7252 N$7254 N$7137 N$7139 "Waveguide Crossing" sch_x=120 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1882 N$7256 N$7258 N$7141 N$7143 "Waveguide Crossing" sch_x=120 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1883 N$7260 N$7262 N$7145 N$7147 "Waveguide Crossing" sch_x=120 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1884 N$7264 N$7266 N$7149 N$7151 "Waveguide Crossing" sch_x=120 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1885 N$7268 N$7270 N$7153 N$7155 "Waveguide Crossing" sch_x=120 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1886 N$7272 N$7274 N$7157 N$7159 "Waveguide Crossing" sch_x=120 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1887 N$7276 N$7278 N$7161 N$7163 "Waveguide Crossing" sch_x=120 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1888 N$7280 N$7282 N$7165 N$7167 "Waveguide Crossing" sch_x=120 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1889 N$7284 N$7286 N$7169 N$7171 "Waveguide Crossing" sch_x=120 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1890 N$7288 N$7290 N$7173 N$7175 "Waveguide Crossing" sch_x=120 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1891 N$7292 N$7294 N$7177 N$7179 "Waveguide Crossing" sch_x=120 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1892 N$7296 N$7298 N$7181 N$7183 "Waveguide Crossing" sch_x=120 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1893 N$7300 N$7302 N$7185 N$7187 "Waveguide Crossing" sch_x=120 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1894 N$7304 N$7306 N$7189 N$7191 "Waveguide Crossing" sch_x=120 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1895 N$7308 N$7310 N$7193 N$7195 "Waveguide Crossing" sch_x=120 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1896 N$7312 N$7314 N$7197 N$7199 "Waveguide Crossing" sch_x=120 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1897 N$7316 N$7318 N$7201 N$7203 "Waveguide Crossing" sch_x=120 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1898 N$7320 N$8951 N$7205 N$7207 "Waveguide Crossing" sch_x=120 sch_y=-28 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1899 N$8839 N$7322 N$7209 N$7211 "Waveguide Crossing" sch_x=118 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1900 N$7324 N$7326 N$7213 N$7215 "Waveguide Crossing" sch_x=118 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1901 N$7328 N$7330 N$7217 N$7219 "Waveguide Crossing" sch_x=118 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1902 N$7332 N$7334 N$7221 N$7223 "Waveguide Crossing" sch_x=118 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1903 N$7336 N$7338 N$7225 N$7227 "Waveguide Crossing" sch_x=118 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1904 N$7340 N$7342 N$7229 N$7231 "Waveguide Crossing" sch_x=118 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1905 N$7344 N$7346 N$7233 N$7235 "Waveguide Crossing" sch_x=118 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1906 N$7348 N$7350 N$7237 N$7239 "Waveguide Crossing" sch_x=118 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1907 N$7352 N$7354 N$7241 N$7243 "Waveguide Crossing" sch_x=118 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1908 N$7356 N$7358 N$7245 N$7247 "Waveguide Crossing" sch_x=118 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1909 N$7360 N$7362 N$7249 N$7251 "Waveguide Crossing" sch_x=118 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1910 N$7364 N$7366 N$7253 N$7255 "Waveguide Crossing" sch_x=118 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1911 N$7368 N$7370 N$7257 N$7259 "Waveguide Crossing" sch_x=118 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1912 N$7372 N$7374 N$7261 N$7263 "Waveguide Crossing" sch_x=118 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1913 N$7376 N$7378 N$7265 N$7267 "Waveguide Crossing" sch_x=118 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1914 N$7380 N$7382 N$7269 N$7271 "Waveguide Crossing" sch_x=118 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1915 N$7384 N$7386 N$7273 N$7275 "Waveguide Crossing" sch_x=118 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1916 N$7388 N$7390 N$7277 N$7279 "Waveguide Crossing" sch_x=118 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1917 N$7392 N$7394 N$7281 N$7283 "Waveguide Crossing" sch_x=118 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1918 N$7396 N$7398 N$7285 N$7287 "Waveguide Crossing" sch_x=118 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1919 N$7400 N$7402 N$7289 N$7291 "Waveguide Crossing" sch_x=118 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1920 N$7404 N$7406 N$7293 N$7295 "Waveguide Crossing" sch_x=118 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1921 N$7408 N$7410 N$7297 N$7299 "Waveguide Crossing" sch_x=118 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1922 N$7412 N$7414 N$7301 N$7303 "Waveguide Crossing" sch_x=118 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1923 N$7416 N$7418 N$7305 N$7307 "Waveguide Crossing" sch_x=118 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1924 N$7420 N$7422 N$7309 N$7311 "Waveguide Crossing" sch_x=118 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1925 N$7424 N$7426 N$7313 N$7315 "Waveguide Crossing" sch_x=118 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1926 N$7428 N$8949 N$7317 N$7319 "Waveguide Crossing" sch_x=118 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1927 N$8841 N$7430 N$7321 N$7323 "Waveguide Crossing" sch_x=116 sch_y=26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1928 N$7432 N$7434 N$7325 N$7327 "Waveguide Crossing" sch_x=116 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1929 N$7436 N$7438 N$7329 N$7331 "Waveguide Crossing" sch_x=116 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1930 N$7440 N$7442 N$7333 N$7335 "Waveguide Crossing" sch_x=116 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1931 N$7444 N$7446 N$7337 N$7339 "Waveguide Crossing" sch_x=116 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1932 N$7448 N$7450 N$7341 N$7343 "Waveguide Crossing" sch_x=116 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1933 N$7452 N$7454 N$7345 N$7347 "Waveguide Crossing" sch_x=116 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1934 N$7456 N$7458 N$7349 N$7351 "Waveguide Crossing" sch_x=116 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1935 N$7460 N$7462 N$7353 N$7355 "Waveguide Crossing" sch_x=116 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1936 N$7464 N$7466 N$7357 N$7359 "Waveguide Crossing" sch_x=116 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1937 N$7468 N$7470 N$7361 N$7363 "Waveguide Crossing" sch_x=116 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1938 N$7472 N$7474 N$7365 N$7367 "Waveguide Crossing" sch_x=116 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1939 N$7476 N$7478 N$7369 N$7371 "Waveguide Crossing" sch_x=116 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1940 N$7480 N$7482 N$7373 N$7375 "Waveguide Crossing" sch_x=116 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1941 N$7484 N$7486 N$7377 N$7379 "Waveguide Crossing" sch_x=116 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1942 N$7488 N$7490 N$7381 N$7383 "Waveguide Crossing" sch_x=116 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1943 N$7492 N$7494 N$7385 N$7387 "Waveguide Crossing" sch_x=116 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1944 N$7496 N$7498 N$7389 N$7391 "Waveguide Crossing" sch_x=116 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1945 N$7500 N$7502 N$7393 N$7395 "Waveguide Crossing" sch_x=116 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1946 N$7504 N$7506 N$7397 N$7399 "Waveguide Crossing" sch_x=116 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1947 N$7508 N$7510 N$7401 N$7403 "Waveguide Crossing" sch_x=116 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1948 N$7512 N$7514 N$7405 N$7407 "Waveguide Crossing" sch_x=116 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1949 N$7516 N$7518 N$7409 N$7411 "Waveguide Crossing" sch_x=116 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1950 N$7520 N$7522 N$7413 N$7415 "Waveguide Crossing" sch_x=116 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1951 N$7524 N$7526 N$7417 N$7419 "Waveguide Crossing" sch_x=116 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1952 N$7528 N$7530 N$7421 N$7423 "Waveguide Crossing" sch_x=116 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1953 N$7532 N$8947 N$7425 N$7427 "Waveguide Crossing" sch_x=116 sch_y=-26 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1954 N$8843 N$7534 N$7429 N$7431 "Waveguide Crossing" sch_x=114 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1955 N$7536 N$7538 N$7433 N$7435 "Waveguide Crossing" sch_x=114 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1956 N$7540 N$7542 N$7437 N$7439 "Waveguide Crossing" sch_x=114 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1957 N$7544 N$7546 N$7441 N$7443 "Waveguide Crossing" sch_x=114 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1958 N$7548 N$7550 N$7445 N$7447 "Waveguide Crossing" sch_x=114 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1959 N$7552 N$7554 N$7449 N$7451 "Waveguide Crossing" sch_x=114 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1960 N$7556 N$7558 N$7453 N$7455 "Waveguide Crossing" sch_x=114 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1961 N$7560 N$7562 N$7457 N$7459 "Waveguide Crossing" sch_x=114 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1962 N$7564 N$7566 N$7461 N$7463 "Waveguide Crossing" sch_x=114 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1963 N$7568 N$7570 N$7465 N$7467 "Waveguide Crossing" sch_x=114 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1964 N$7572 N$7574 N$7469 N$7471 "Waveguide Crossing" sch_x=114 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1965 N$7576 N$7578 N$7473 N$7475 "Waveguide Crossing" sch_x=114 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1966 N$7580 N$7582 N$7477 N$7479 "Waveguide Crossing" sch_x=114 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1967 N$7584 N$7586 N$7481 N$7483 "Waveguide Crossing" sch_x=114 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1968 N$7588 N$7590 N$7485 N$7487 "Waveguide Crossing" sch_x=114 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1969 N$7592 N$7594 N$7489 N$7491 "Waveguide Crossing" sch_x=114 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1970 N$7596 N$7598 N$7493 N$7495 "Waveguide Crossing" sch_x=114 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1971 N$7600 N$7602 N$7497 N$7499 "Waveguide Crossing" sch_x=114 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1972 N$7604 N$7606 N$7501 N$7503 "Waveguide Crossing" sch_x=114 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1973 N$7608 N$7610 N$7505 N$7507 "Waveguide Crossing" sch_x=114 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1974 N$7612 N$7614 N$7509 N$7511 "Waveguide Crossing" sch_x=114 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1975 N$7616 N$7618 N$7513 N$7515 "Waveguide Crossing" sch_x=114 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1976 N$7620 N$7622 N$7517 N$7519 "Waveguide Crossing" sch_x=114 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1977 N$7624 N$7626 N$7521 N$7523 "Waveguide Crossing" sch_x=114 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1978 N$7628 N$7630 N$7525 N$7527 "Waveguide Crossing" sch_x=114 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1979 N$7632 N$8945 N$7529 N$7531 "Waveguide Crossing" sch_x=114 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1980 N$8845 N$7634 N$7533 N$7535 "Waveguide Crossing" sch_x=112 sch_y=24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1981 N$7636 N$7638 N$7537 N$7539 "Waveguide Crossing" sch_x=112 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1982 N$7640 N$7642 N$7541 N$7543 "Waveguide Crossing" sch_x=112 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1983 N$7644 N$7646 N$7545 N$7547 "Waveguide Crossing" sch_x=112 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1984 N$7648 N$7650 N$7549 N$7551 "Waveguide Crossing" sch_x=112 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1985 N$7652 N$7654 N$7553 N$7555 "Waveguide Crossing" sch_x=112 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1986 N$7656 N$7658 N$7557 N$7559 "Waveguide Crossing" sch_x=112 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1987 N$7660 N$7662 N$7561 N$7563 "Waveguide Crossing" sch_x=112 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1988 N$7664 N$7666 N$7565 N$7567 "Waveguide Crossing" sch_x=112 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1989 N$7668 N$7670 N$7569 N$7571 "Waveguide Crossing" sch_x=112 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1990 N$7672 N$7674 N$7573 N$7575 "Waveguide Crossing" sch_x=112 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1991 N$7676 N$7678 N$7577 N$7579 "Waveguide Crossing" sch_x=112 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1992 N$7680 N$7682 N$7581 N$7583 "Waveguide Crossing" sch_x=112 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1993 N$7684 N$7686 N$7585 N$7587 "Waveguide Crossing" sch_x=112 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1994 N$7688 N$7690 N$7589 N$7591 "Waveguide Crossing" sch_x=112 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1995 N$7692 N$7694 N$7593 N$7595 "Waveguide Crossing" sch_x=112 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1996 N$7696 N$7698 N$7597 N$7599 "Waveguide Crossing" sch_x=112 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1997 N$7700 N$7702 N$7601 N$7603 "Waveguide Crossing" sch_x=112 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1998 N$7704 N$7706 N$7605 N$7607 "Waveguide Crossing" sch_x=112 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C1999 N$7708 N$7710 N$7609 N$7611 "Waveguide Crossing" sch_x=112 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2000 N$7712 N$7714 N$7613 N$7615 "Waveguide Crossing" sch_x=112 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2001 N$7716 N$7718 N$7617 N$7619 "Waveguide Crossing" sch_x=112 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2002 N$7720 N$7722 N$7621 N$7623 "Waveguide Crossing" sch_x=112 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2003 N$7724 N$7726 N$7625 N$7627 "Waveguide Crossing" sch_x=112 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2004 N$7728 N$8943 N$7629 N$7631 "Waveguide Crossing" sch_x=112 sch_y=-24 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2005 N$8847 N$7730 N$7633 N$7635 "Waveguide Crossing" sch_x=110 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2006 N$7732 N$7734 N$7637 N$7639 "Waveguide Crossing" sch_x=110 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2007 N$7736 N$7738 N$7641 N$7643 "Waveguide Crossing" sch_x=110 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2008 N$7740 N$7742 N$7645 N$7647 "Waveguide Crossing" sch_x=110 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2009 N$7744 N$7746 N$7649 N$7651 "Waveguide Crossing" sch_x=110 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2010 N$7748 N$7750 N$7653 N$7655 "Waveguide Crossing" sch_x=110 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2011 N$7752 N$7754 N$7657 N$7659 "Waveguide Crossing" sch_x=110 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2012 N$7756 N$7758 N$7661 N$7663 "Waveguide Crossing" sch_x=110 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2013 N$7760 N$7762 N$7665 N$7667 "Waveguide Crossing" sch_x=110 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2014 N$7764 N$7766 N$7669 N$7671 "Waveguide Crossing" sch_x=110 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2015 N$7768 N$7770 N$7673 N$7675 "Waveguide Crossing" sch_x=110 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2016 N$7772 N$7774 N$7677 N$7679 "Waveguide Crossing" sch_x=110 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2017 N$7776 N$7778 N$7681 N$7683 "Waveguide Crossing" sch_x=110 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2018 N$7780 N$7782 N$7685 N$7687 "Waveguide Crossing" sch_x=110 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2019 N$7784 N$7786 N$7689 N$7691 "Waveguide Crossing" sch_x=110 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2020 N$7788 N$7790 N$7693 N$7695 "Waveguide Crossing" sch_x=110 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2021 N$7792 N$7794 N$7697 N$7699 "Waveguide Crossing" sch_x=110 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2022 N$7796 N$7798 N$7701 N$7703 "Waveguide Crossing" sch_x=110 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2023 N$7800 N$7802 N$7705 N$7707 "Waveguide Crossing" sch_x=110 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2024 N$7804 N$7806 N$7709 N$7711 "Waveguide Crossing" sch_x=110 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2025 N$7808 N$7810 N$7713 N$7715 "Waveguide Crossing" sch_x=110 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2026 N$7812 N$7814 N$7717 N$7719 "Waveguide Crossing" sch_x=110 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2027 N$7816 N$7818 N$7721 N$7723 "Waveguide Crossing" sch_x=110 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2028 N$7820 N$8941 N$7725 N$7727 "Waveguide Crossing" sch_x=110 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2029 N$8849 N$7822 N$7729 N$7731 "Waveguide Crossing" sch_x=108 sch_y=22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2030 N$7824 N$7826 N$7733 N$7735 "Waveguide Crossing" sch_x=108 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2031 N$7828 N$7830 N$7737 N$7739 "Waveguide Crossing" sch_x=108 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2032 N$7832 N$7834 N$7741 N$7743 "Waveguide Crossing" sch_x=108 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2033 N$7836 N$7838 N$7745 N$7747 "Waveguide Crossing" sch_x=108 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2034 N$7840 N$7842 N$7749 N$7751 "Waveguide Crossing" sch_x=108 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2035 N$7844 N$7846 N$7753 N$7755 "Waveguide Crossing" sch_x=108 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2036 N$7848 N$7850 N$7757 N$7759 "Waveguide Crossing" sch_x=108 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2037 N$7852 N$7854 N$7761 N$7763 "Waveguide Crossing" sch_x=108 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2038 N$7856 N$7858 N$7765 N$7767 "Waveguide Crossing" sch_x=108 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2039 N$7860 N$7862 N$7769 N$7771 "Waveguide Crossing" sch_x=108 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2040 N$7864 N$7866 N$7773 N$7775 "Waveguide Crossing" sch_x=108 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2041 N$7868 N$7870 N$7777 N$7779 "Waveguide Crossing" sch_x=108 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2042 N$7872 N$7874 N$7781 N$7783 "Waveguide Crossing" sch_x=108 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2043 N$7876 N$7878 N$7785 N$7787 "Waveguide Crossing" sch_x=108 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2044 N$7880 N$7882 N$7789 N$7791 "Waveguide Crossing" sch_x=108 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2045 N$7884 N$7886 N$7793 N$7795 "Waveguide Crossing" sch_x=108 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2046 N$7888 N$7890 N$7797 N$7799 "Waveguide Crossing" sch_x=108 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2047 N$7892 N$7894 N$7801 N$7803 "Waveguide Crossing" sch_x=108 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2048 N$7896 N$7898 N$7805 N$7807 "Waveguide Crossing" sch_x=108 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2049 N$7900 N$7902 N$7809 N$7811 "Waveguide Crossing" sch_x=108 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2050 N$7904 N$7906 N$7813 N$7815 "Waveguide Crossing" sch_x=108 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2051 N$7908 N$8939 N$7817 N$7819 "Waveguide Crossing" sch_x=108 sch_y=-22 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2052 N$8851 N$7910 N$7821 N$7823 "Waveguide Crossing" sch_x=106 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2053 N$7912 N$7914 N$7825 N$7827 "Waveguide Crossing" sch_x=106 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2054 N$7916 N$7918 N$7829 N$7831 "Waveguide Crossing" sch_x=106 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2055 N$7920 N$7922 N$7833 N$7835 "Waveguide Crossing" sch_x=106 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2056 N$7924 N$7926 N$7837 N$7839 "Waveguide Crossing" sch_x=106 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2057 N$7928 N$7930 N$7841 N$7843 "Waveguide Crossing" sch_x=106 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2058 N$7932 N$7934 N$7845 N$7847 "Waveguide Crossing" sch_x=106 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2059 N$7936 N$7938 N$7849 N$7851 "Waveguide Crossing" sch_x=106 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2060 N$7940 N$7942 N$7853 N$7855 "Waveguide Crossing" sch_x=106 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2061 N$7944 N$7946 N$7857 N$7859 "Waveguide Crossing" sch_x=106 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2062 N$7948 N$7950 N$7861 N$7863 "Waveguide Crossing" sch_x=106 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2063 N$7952 N$7954 N$7865 N$7867 "Waveguide Crossing" sch_x=106 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2064 N$7956 N$7958 N$7869 N$7871 "Waveguide Crossing" sch_x=106 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2065 N$7960 N$7962 N$7873 N$7875 "Waveguide Crossing" sch_x=106 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2066 N$7964 N$7966 N$7877 N$7879 "Waveguide Crossing" sch_x=106 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2067 N$7968 N$7970 N$7881 N$7883 "Waveguide Crossing" sch_x=106 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2068 N$7972 N$7974 N$7885 N$7887 "Waveguide Crossing" sch_x=106 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2069 N$7976 N$7978 N$7889 N$7891 "Waveguide Crossing" sch_x=106 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2070 N$7980 N$7982 N$7893 N$7895 "Waveguide Crossing" sch_x=106 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2071 N$7984 N$7986 N$7897 N$7899 "Waveguide Crossing" sch_x=106 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2072 N$7988 N$7990 N$7901 N$7903 "Waveguide Crossing" sch_x=106 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2073 N$7992 N$8937 N$7905 N$7907 "Waveguide Crossing" sch_x=106 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2074 N$8853 N$7994 N$7909 N$7911 "Waveguide Crossing" sch_x=104 sch_y=20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2075 N$7996 N$7998 N$7913 N$7915 "Waveguide Crossing" sch_x=104 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2076 N$8000 N$8002 N$7917 N$7919 "Waveguide Crossing" sch_x=104 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2077 N$8004 N$8006 N$7921 N$7923 "Waveguide Crossing" sch_x=104 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2078 N$8008 N$8010 N$7925 N$7927 "Waveguide Crossing" sch_x=104 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2079 N$8012 N$8014 N$7929 N$7931 "Waveguide Crossing" sch_x=104 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2080 N$8016 N$8018 N$7933 N$7935 "Waveguide Crossing" sch_x=104 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2081 N$8020 N$8022 N$7937 N$7939 "Waveguide Crossing" sch_x=104 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2082 N$8024 N$8026 N$7941 N$7943 "Waveguide Crossing" sch_x=104 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2083 N$8028 N$8030 N$7945 N$7947 "Waveguide Crossing" sch_x=104 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2084 N$8032 N$8034 N$7949 N$7951 "Waveguide Crossing" sch_x=104 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2085 N$8036 N$8038 N$7953 N$7955 "Waveguide Crossing" sch_x=104 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2086 N$8040 N$8042 N$7957 N$7959 "Waveguide Crossing" sch_x=104 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2087 N$8044 N$8046 N$7961 N$7963 "Waveguide Crossing" sch_x=104 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2088 N$8048 N$8050 N$7965 N$7967 "Waveguide Crossing" sch_x=104 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2089 N$8052 N$8054 N$7969 N$7971 "Waveguide Crossing" sch_x=104 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2090 N$8056 N$8058 N$7973 N$7975 "Waveguide Crossing" sch_x=104 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2091 N$8060 N$8062 N$7977 N$7979 "Waveguide Crossing" sch_x=104 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2092 N$8064 N$8066 N$7981 N$7983 "Waveguide Crossing" sch_x=104 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2093 N$8068 N$8070 N$7985 N$7987 "Waveguide Crossing" sch_x=104 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2094 N$8072 N$8935 N$7989 N$7991 "Waveguide Crossing" sch_x=104 sch_y=-20 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2095 N$8855 N$8074 N$7993 N$7995 "Waveguide Crossing" sch_x=102 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2096 N$8076 N$8078 N$7997 N$7999 "Waveguide Crossing" sch_x=102 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2097 N$8080 N$8082 N$8001 N$8003 "Waveguide Crossing" sch_x=102 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2098 N$8084 N$8086 N$8005 N$8007 "Waveguide Crossing" sch_x=102 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2099 N$8088 N$8090 N$8009 N$8011 "Waveguide Crossing" sch_x=102 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2100 N$8092 N$8094 N$8013 N$8015 "Waveguide Crossing" sch_x=102 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2101 N$8096 N$8098 N$8017 N$8019 "Waveguide Crossing" sch_x=102 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2102 N$8100 N$8102 N$8021 N$8023 "Waveguide Crossing" sch_x=102 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2103 N$8104 N$8106 N$8025 N$8027 "Waveguide Crossing" sch_x=102 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2104 N$8108 N$8110 N$8029 N$8031 "Waveguide Crossing" sch_x=102 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2105 N$8112 N$8114 N$8033 N$8035 "Waveguide Crossing" sch_x=102 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2106 N$8116 N$8118 N$8037 N$8039 "Waveguide Crossing" sch_x=102 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2107 N$8120 N$8122 N$8041 N$8043 "Waveguide Crossing" sch_x=102 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2108 N$8124 N$8126 N$8045 N$8047 "Waveguide Crossing" sch_x=102 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2109 N$8128 N$8130 N$8049 N$8051 "Waveguide Crossing" sch_x=102 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2110 N$8132 N$8134 N$8053 N$8055 "Waveguide Crossing" sch_x=102 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2111 N$8136 N$8138 N$8057 N$8059 "Waveguide Crossing" sch_x=102 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2112 N$8140 N$8142 N$8061 N$8063 "Waveguide Crossing" sch_x=102 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2113 N$8144 N$8146 N$8065 N$8067 "Waveguide Crossing" sch_x=102 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2114 N$8148 N$8933 N$8069 N$8071 "Waveguide Crossing" sch_x=102 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2115 N$8857 N$8150 N$8073 N$8075 "Waveguide Crossing" sch_x=100 sch_y=18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2116 N$8152 N$8154 N$8077 N$8079 "Waveguide Crossing" sch_x=100 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2117 N$8156 N$8158 N$8081 N$8083 "Waveguide Crossing" sch_x=100 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2118 N$8160 N$8162 N$8085 N$8087 "Waveguide Crossing" sch_x=100 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2119 N$8164 N$8166 N$8089 N$8091 "Waveguide Crossing" sch_x=100 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2120 N$8168 N$8170 N$8093 N$8095 "Waveguide Crossing" sch_x=100 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2121 N$8172 N$8174 N$8097 N$8099 "Waveguide Crossing" sch_x=100 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2122 N$8176 N$8178 N$8101 N$8103 "Waveguide Crossing" sch_x=100 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2123 N$8180 N$8182 N$8105 N$8107 "Waveguide Crossing" sch_x=100 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2124 N$8184 N$8186 N$8109 N$8111 "Waveguide Crossing" sch_x=100 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2125 N$8188 N$8190 N$8113 N$8115 "Waveguide Crossing" sch_x=100 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2126 N$8192 N$8194 N$8117 N$8119 "Waveguide Crossing" sch_x=100 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2127 N$8196 N$8198 N$8121 N$8123 "Waveguide Crossing" sch_x=100 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2128 N$8200 N$8202 N$8125 N$8127 "Waveguide Crossing" sch_x=100 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2129 N$8204 N$8206 N$8129 N$8131 "Waveguide Crossing" sch_x=100 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2130 N$8208 N$8210 N$8133 N$8135 "Waveguide Crossing" sch_x=100 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2131 N$8212 N$8214 N$8137 N$8139 "Waveguide Crossing" sch_x=100 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2132 N$8216 N$8218 N$8141 N$8143 "Waveguide Crossing" sch_x=100 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2133 N$8220 N$8931 N$8145 N$8147 "Waveguide Crossing" sch_x=100 sch_y=-18 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2134 N$8859 N$8222 N$8149 N$8151 "Waveguide Crossing" sch_x=98 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2135 N$8224 N$8226 N$8153 N$8155 "Waveguide Crossing" sch_x=98 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2136 N$8228 N$8230 N$8157 N$8159 "Waveguide Crossing" sch_x=98 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2137 N$8232 N$8234 N$8161 N$8163 "Waveguide Crossing" sch_x=98 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2138 N$8236 N$8238 N$8165 N$8167 "Waveguide Crossing" sch_x=98 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2139 N$8240 N$8242 N$8169 N$8171 "Waveguide Crossing" sch_x=98 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2140 N$8244 N$8246 N$8173 N$8175 "Waveguide Crossing" sch_x=98 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2141 N$8248 N$8250 N$8177 N$8179 "Waveguide Crossing" sch_x=98 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2142 N$8252 N$8254 N$8181 N$8183 "Waveguide Crossing" sch_x=98 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2143 N$8256 N$8258 N$8185 N$8187 "Waveguide Crossing" sch_x=98 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2144 N$8260 N$8262 N$8189 N$8191 "Waveguide Crossing" sch_x=98 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2145 N$8264 N$8266 N$8193 N$8195 "Waveguide Crossing" sch_x=98 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2146 N$8268 N$8270 N$8197 N$8199 "Waveguide Crossing" sch_x=98 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2147 N$8272 N$8274 N$8201 N$8203 "Waveguide Crossing" sch_x=98 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2148 N$8276 N$8278 N$8205 N$8207 "Waveguide Crossing" sch_x=98 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2149 N$8280 N$8282 N$8209 N$8211 "Waveguide Crossing" sch_x=98 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2150 N$8284 N$8286 N$8213 N$8215 "Waveguide Crossing" sch_x=98 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2151 N$8288 N$8929 N$8217 N$8219 "Waveguide Crossing" sch_x=98 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2152 N$8861 N$8290 N$8221 N$8223 "Waveguide Crossing" sch_x=96 sch_y=16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2153 N$8292 N$8294 N$8225 N$8227 "Waveguide Crossing" sch_x=96 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2154 N$8296 N$8298 N$8229 N$8231 "Waveguide Crossing" sch_x=96 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2155 N$8300 N$8302 N$8233 N$8235 "Waveguide Crossing" sch_x=96 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2156 N$8304 N$8306 N$8237 N$8239 "Waveguide Crossing" sch_x=96 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2157 N$8308 N$8310 N$8241 N$8243 "Waveguide Crossing" sch_x=96 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2158 N$8312 N$8314 N$8245 N$8247 "Waveguide Crossing" sch_x=96 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2159 N$8316 N$8318 N$8249 N$8251 "Waveguide Crossing" sch_x=96 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2160 N$8320 N$8322 N$8253 N$8255 "Waveguide Crossing" sch_x=96 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2161 N$8324 N$8326 N$8257 N$8259 "Waveguide Crossing" sch_x=96 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2162 N$8328 N$8330 N$8261 N$8263 "Waveguide Crossing" sch_x=96 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2163 N$8332 N$8334 N$8265 N$8267 "Waveguide Crossing" sch_x=96 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2164 N$8336 N$8338 N$8269 N$8271 "Waveguide Crossing" sch_x=96 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2165 N$8340 N$8342 N$8273 N$8275 "Waveguide Crossing" sch_x=96 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2166 N$8344 N$8346 N$8277 N$8279 "Waveguide Crossing" sch_x=96 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2167 N$8348 N$8350 N$8281 N$8283 "Waveguide Crossing" sch_x=96 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2168 N$8352 N$8927 N$8285 N$8287 "Waveguide Crossing" sch_x=96 sch_y=-16 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2169 N$8863 N$8354 N$8289 N$8291 "Waveguide Crossing" sch_x=94 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2170 N$8356 N$8358 N$8293 N$8295 "Waveguide Crossing" sch_x=94 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2171 N$8360 N$8362 N$8297 N$8299 "Waveguide Crossing" sch_x=94 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2172 N$8364 N$8366 N$8301 N$8303 "Waveguide Crossing" sch_x=94 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2173 N$8368 N$8370 N$8305 N$8307 "Waveguide Crossing" sch_x=94 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2174 N$8372 N$8374 N$8309 N$8311 "Waveguide Crossing" sch_x=94 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2175 N$8376 N$8378 N$8313 N$8315 "Waveguide Crossing" sch_x=94 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2176 N$8380 N$8382 N$8317 N$8319 "Waveguide Crossing" sch_x=94 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2177 N$8384 N$8386 N$8321 N$8323 "Waveguide Crossing" sch_x=94 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2178 N$8388 N$8390 N$8325 N$8327 "Waveguide Crossing" sch_x=94 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2179 N$8392 N$8394 N$8329 N$8331 "Waveguide Crossing" sch_x=94 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2180 N$8396 N$8398 N$8333 N$8335 "Waveguide Crossing" sch_x=94 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2181 N$8400 N$8402 N$8337 N$8339 "Waveguide Crossing" sch_x=94 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2182 N$8404 N$8406 N$8341 N$8343 "Waveguide Crossing" sch_x=94 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2183 N$8408 N$8410 N$8345 N$8347 "Waveguide Crossing" sch_x=94 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2184 N$8412 N$8925 N$8349 N$8351 "Waveguide Crossing" sch_x=94 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2185 N$8865 N$8414 N$8353 N$8355 "Waveguide Crossing" sch_x=92 sch_y=14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2186 N$8416 N$8418 N$8357 N$8359 "Waveguide Crossing" sch_x=92 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2187 N$8420 N$8422 N$8361 N$8363 "Waveguide Crossing" sch_x=92 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2188 N$8424 N$8426 N$8365 N$8367 "Waveguide Crossing" sch_x=92 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2189 N$8428 N$8430 N$8369 N$8371 "Waveguide Crossing" sch_x=92 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2190 N$8432 N$8434 N$8373 N$8375 "Waveguide Crossing" sch_x=92 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2191 N$8436 N$8438 N$8377 N$8379 "Waveguide Crossing" sch_x=92 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2192 N$8440 N$8442 N$8381 N$8383 "Waveguide Crossing" sch_x=92 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2193 N$8444 N$8446 N$8385 N$8387 "Waveguide Crossing" sch_x=92 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2194 N$8448 N$8450 N$8389 N$8391 "Waveguide Crossing" sch_x=92 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2195 N$8452 N$8454 N$8393 N$8395 "Waveguide Crossing" sch_x=92 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2196 N$8456 N$8458 N$8397 N$8399 "Waveguide Crossing" sch_x=92 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2197 N$8460 N$8462 N$8401 N$8403 "Waveguide Crossing" sch_x=92 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2198 N$8464 N$8466 N$8405 N$8407 "Waveguide Crossing" sch_x=92 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2199 N$8468 N$8923 N$8409 N$8411 "Waveguide Crossing" sch_x=92 sch_y=-14 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2200 N$8867 N$8470 N$8413 N$8415 "Waveguide Crossing" sch_x=90 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2201 N$8472 N$8474 N$8417 N$8419 "Waveguide Crossing" sch_x=90 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2202 N$8476 N$8478 N$8421 N$8423 "Waveguide Crossing" sch_x=90 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2203 N$8480 N$8482 N$8425 N$8427 "Waveguide Crossing" sch_x=90 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2204 N$8484 N$8486 N$8429 N$8431 "Waveguide Crossing" sch_x=90 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2205 N$8488 N$8490 N$8433 N$8435 "Waveguide Crossing" sch_x=90 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2206 N$8492 N$8494 N$8437 N$8439 "Waveguide Crossing" sch_x=90 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2207 N$8496 N$8498 N$8441 N$8443 "Waveguide Crossing" sch_x=90 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2208 N$8500 N$8502 N$8445 N$8447 "Waveguide Crossing" sch_x=90 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2209 N$8504 N$8506 N$8449 N$8451 "Waveguide Crossing" sch_x=90 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2210 N$8508 N$8510 N$8453 N$8455 "Waveguide Crossing" sch_x=90 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2211 N$8512 N$8514 N$8457 N$8459 "Waveguide Crossing" sch_x=90 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2212 N$8516 N$8518 N$8461 N$8463 "Waveguide Crossing" sch_x=90 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2213 N$8520 N$8921 N$8465 N$8467 "Waveguide Crossing" sch_x=90 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2214 N$8869 N$8522 N$8469 N$8471 "Waveguide Crossing" sch_x=88 sch_y=12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2215 N$8524 N$8526 N$8473 N$8475 "Waveguide Crossing" sch_x=88 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2216 N$8528 N$8530 N$8477 N$8479 "Waveguide Crossing" sch_x=88 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2217 N$8532 N$8534 N$8481 N$8483 "Waveguide Crossing" sch_x=88 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2218 N$8536 N$8538 N$8485 N$8487 "Waveguide Crossing" sch_x=88 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2219 N$8540 N$8542 N$8489 N$8491 "Waveguide Crossing" sch_x=88 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2220 N$8544 N$8546 N$8493 N$8495 "Waveguide Crossing" sch_x=88 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2221 N$8548 N$8550 N$8497 N$8499 "Waveguide Crossing" sch_x=88 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2222 N$8552 N$8554 N$8501 N$8503 "Waveguide Crossing" sch_x=88 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2223 N$8556 N$8558 N$8505 N$8507 "Waveguide Crossing" sch_x=88 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2224 N$8560 N$8562 N$8509 N$8511 "Waveguide Crossing" sch_x=88 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2225 N$8564 N$8566 N$8513 N$8515 "Waveguide Crossing" sch_x=88 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2226 N$8568 N$8919 N$8517 N$8519 "Waveguide Crossing" sch_x=88 sch_y=-12 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2227 N$8871 N$8570 N$8521 N$8523 "Waveguide Crossing" sch_x=86 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2228 N$8572 N$8574 N$8525 N$8527 "Waveguide Crossing" sch_x=86 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2229 N$8576 N$8578 N$8529 N$8531 "Waveguide Crossing" sch_x=86 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2230 N$8580 N$8582 N$8533 N$8535 "Waveguide Crossing" sch_x=86 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2231 N$8584 N$8586 N$8537 N$8539 "Waveguide Crossing" sch_x=86 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2232 N$8588 N$8590 N$8541 N$8543 "Waveguide Crossing" sch_x=86 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2233 N$8592 N$8594 N$8545 N$8547 "Waveguide Crossing" sch_x=86 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2234 N$8596 N$8598 N$8549 N$8551 "Waveguide Crossing" sch_x=86 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2235 N$8600 N$8602 N$8553 N$8555 "Waveguide Crossing" sch_x=86 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2236 N$8604 N$8606 N$8557 N$8559 "Waveguide Crossing" sch_x=86 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2237 N$8608 N$8610 N$8561 N$8563 "Waveguide Crossing" sch_x=86 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2238 N$8612 N$8917 N$8565 N$8567 "Waveguide Crossing" sch_x=86 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2239 N$8873 N$8614 N$8569 N$8571 "Waveguide Crossing" sch_x=84 sch_y=10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2240 N$8616 N$8618 N$8573 N$8575 "Waveguide Crossing" sch_x=84 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2241 N$8620 N$8622 N$8577 N$8579 "Waveguide Crossing" sch_x=84 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2242 N$8624 N$8626 N$8581 N$8583 "Waveguide Crossing" sch_x=84 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2243 N$8628 N$8630 N$8585 N$8587 "Waveguide Crossing" sch_x=84 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2244 N$8632 N$8634 N$8589 N$8591 "Waveguide Crossing" sch_x=84 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2245 N$8636 N$8638 N$8593 N$8595 "Waveguide Crossing" sch_x=84 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2246 N$8640 N$8642 N$8597 N$8599 "Waveguide Crossing" sch_x=84 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2247 N$8644 N$8646 N$8601 N$8603 "Waveguide Crossing" sch_x=84 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2248 N$8648 N$8650 N$8605 N$8607 "Waveguide Crossing" sch_x=84 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2249 N$8652 N$8915 N$8609 N$8611 "Waveguide Crossing" sch_x=84 sch_y=-10 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2250 N$8875 N$8654 N$8613 N$8615 "Waveguide Crossing" sch_x=82 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2251 N$8656 N$8658 N$8617 N$8619 "Waveguide Crossing" sch_x=82 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2252 N$8660 N$8662 N$8621 N$8623 "Waveguide Crossing" sch_x=82 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2253 N$8664 N$8666 N$8625 N$8627 "Waveguide Crossing" sch_x=82 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2254 N$8668 N$8670 N$8629 N$8631 "Waveguide Crossing" sch_x=82 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2255 N$8672 N$8674 N$8633 N$8635 "Waveguide Crossing" sch_x=82 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2256 N$8676 N$8678 N$8637 N$8639 "Waveguide Crossing" sch_x=82 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2257 N$8680 N$8682 N$8641 N$8643 "Waveguide Crossing" sch_x=82 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2258 N$8684 N$8686 N$8645 N$8647 "Waveguide Crossing" sch_x=82 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2259 N$8688 N$8913 N$8649 N$8651 "Waveguide Crossing" sch_x=82 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2260 N$8877 N$8690 N$8653 N$8655 "Waveguide Crossing" sch_x=80 sch_y=8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2261 N$8692 N$8694 N$8657 N$8659 "Waveguide Crossing" sch_x=80 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2262 N$8696 N$8698 N$8661 N$8663 "Waveguide Crossing" sch_x=80 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2263 N$8700 N$8702 N$8665 N$8667 "Waveguide Crossing" sch_x=80 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2264 N$8704 N$8706 N$8669 N$8671 "Waveguide Crossing" sch_x=80 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2265 N$8708 N$8710 N$8673 N$8675 "Waveguide Crossing" sch_x=80 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2266 N$8712 N$8714 N$8677 N$8679 "Waveguide Crossing" sch_x=80 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2267 N$8716 N$8718 N$8681 N$8683 "Waveguide Crossing" sch_x=80 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2268 N$8720 N$8911 N$8685 N$8687 "Waveguide Crossing" sch_x=80 sch_y=-8 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2269 N$8879 N$8722 N$8689 N$8691 "Waveguide Crossing" sch_x=78 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2270 N$8724 N$8726 N$8693 N$8695 "Waveguide Crossing" sch_x=78 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2271 N$8728 N$8730 N$8697 N$8699 "Waveguide Crossing" sch_x=78 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2272 N$8732 N$8734 N$8701 N$8703 "Waveguide Crossing" sch_x=78 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2273 N$8736 N$8738 N$8705 N$8707 "Waveguide Crossing" sch_x=78 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2274 N$8740 N$8742 N$8709 N$8711 "Waveguide Crossing" sch_x=78 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2275 N$8744 N$8746 N$8713 N$8715 "Waveguide Crossing" sch_x=78 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2276 N$8748 N$8909 N$8717 N$8719 "Waveguide Crossing" sch_x=78 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2277 N$8881 N$8750 N$8721 N$8723 "Waveguide Crossing" sch_x=76 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2278 N$8752 N$8754 N$8725 N$8727 "Waveguide Crossing" sch_x=76 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2279 N$8756 N$8758 N$8729 N$8731 "Waveguide Crossing" sch_x=76 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2280 N$8760 N$8762 N$8733 N$8735 "Waveguide Crossing" sch_x=76 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2281 N$8764 N$8766 N$8737 N$8739 "Waveguide Crossing" sch_x=76 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2282 N$8768 N$8770 N$8741 N$8743 "Waveguide Crossing" sch_x=76 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2283 N$8772 N$8907 N$8745 N$8747 "Waveguide Crossing" sch_x=76 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2284 N$8883 N$8774 N$8749 N$8751 "Waveguide Crossing" sch_x=74 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2285 N$8776 N$8778 N$8753 N$8755 "Waveguide Crossing" sch_x=74 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2286 N$8780 N$8782 N$8757 N$8759 "Waveguide Crossing" sch_x=74 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2287 N$8784 N$8786 N$8761 N$8763 "Waveguide Crossing" sch_x=74 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2288 N$8788 N$8790 N$8765 N$8767 "Waveguide Crossing" sch_x=74 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2289 N$8792 N$8905 N$8769 N$8771 "Waveguide Crossing" sch_x=74 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2290 N$8885 N$8794 N$8773 N$8775 "Waveguide Crossing" sch_x=72 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2291 N$8796 N$8798 N$8777 N$8779 "Waveguide Crossing" sch_x=72 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2292 N$8800 N$8802 N$8781 N$8783 "Waveguide Crossing" sch_x=72 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2293 N$8804 N$8806 N$8785 N$8787 "Waveguide Crossing" sch_x=72 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2294 N$8808 N$8903 N$8789 N$8791 "Waveguide Crossing" sch_x=72 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2295 N$8887 N$8810 N$8793 N$8795 "Waveguide Crossing" sch_x=70 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2296 N$8812 N$8814 N$8797 N$8799 "Waveguide Crossing" sch_x=70 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2297 N$8816 N$8818 N$8801 N$8803 "Waveguide Crossing" sch_x=70 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2298 N$8820 N$8901 N$8805 N$8807 "Waveguide Crossing" sch_x=70 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2299 N$8889 N$8822 N$8809 N$8811 "Waveguide Crossing" sch_x=68 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2300 N$8824 N$8826 N$8813 N$8815 "Waveguide Crossing" sch_x=68 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2301 N$8828 N$8899 N$8817 N$8819 "Waveguide Crossing" sch_x=68 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2302 N$8891 N$8830 N$8821 N$8823 "Waveguide Crossing" sch_x=66 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2303 N$8832 N$8897 N$8825 N$8827 "Waveguide Crossing" sch_x=66 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C2304 N$8893 N$8895 N$8829 N$8831 "Waveguide Crossing" sch_x=64 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1777 N$8957 N$6850 N$9153 N$9154 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1778 N$6852 N$6854 N$9155 N$9156 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1779 N$6856 N$6858 N$9157 N$9158 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1780 N$6860 N$6862 N$9159 N$9160 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1781 N$6864 N$6866 N$9161 N$9162 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1782 N$6868 N$6870 N$9163 N$9164 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1783 N$6872 N$6874 N$9165 N$9166 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1784 N$6876 N$6878 N$9167 N$9168 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1785 N$6880 N$6882 N$9169 N$9170 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1786 N$6884 N$6886 N$9171 N$9172 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1787 N$6888 N$6890 N$9173 N$9174 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1788 N$6892 N$6894 N$9175 N$9176 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1789 N$6896 N$6898 N$9177 N$9178 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1790 N$6900 N$6902 N$9179 N$9180 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1791 N$6904 N$6906 N$9181 N$9182 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1792 N$6908 N$6910 N$9183 N$9184 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1793 N$6912 N$6914 N$9185 N$9186 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1794 N$6916 N$6918 N$9187 N$9188 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1795 N$6920 N$6922 N$9189 N$9190 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1796 N$6924 N$6926 N$9191 N$9192 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1797 N$6928 N$6930 N$9193 N$9194 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1798 N$6932 N$6934 N$9195 N$9196 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1799 N$6936 N$6938 N$9197 N$9198 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1800 N$6940 N$6942 N$9199 N$9200 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1801 N$6944 N$6946 N$9201 N$9202 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1802 N$6948 N$6950 N$9203 N$9204 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1803 N$6952 N$6954 N$9205 N$9206 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1804 N$6956 N$6958 N$9207 N$9208 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1805 N$6960 N$6962 N$9209 N$9210 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1806 N$6964 N$6966 N$9211 N$9212 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1807 N$6968 N$6970 N$9213 N$9214 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1808 N$6972 N$8959 N$9215 N$9216 MMI_switch_ideal library="Design kits/capstone" sch_x=126 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1 N$1 N$2 "Straight Waveguide" sch_x=-4 sch_y=31.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2 N$3 N$4 "Straight Waveguide" sch_x=-5 sch_y=30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3 N$5 N$6 "Straight Waveguide" sch_x=-5 sch_y=29.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4 N$7 N$8 "Straight Waveguide" sch_x=-3 sch_y=30.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W5 N$9 N$10 "Straight Waveguide" sch_x=-3 sch_y=29.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W6 N$11 N$12 "Straight Waveguide" sch_x=-4 sch_y=28.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W7 N$13 N$14 "Straight Waveguide" sch_x=0 sch_y=31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W8 N$15 N$16 "Straight Waveguide" sch_x=-1 sch_y=31.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W9 N$17 N$18 "Straight Waveguide" sch_x=-1 sch_y=30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W10 N$19 N$20 "Straight Waveguide" sch_x=1 sch_y=30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W11 N$21 N$22 "Straight Waveguide" sch_x=1 sch_y=31.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W12 N$23 N$24 "Straight Waveguide" sch_x=0 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W13 N$25 N$26 "Straight Waveguide" sch_x=0 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W14 N$27 N$28 "Straight Waveguide" sch_x=-1 sch_y=29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W15 N$29 N$30 "Straight Waveguide" sch_x=-1 sch_y=28.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W16 N$31 N$32 "Straight Waveguide" sch_x=1 sch_y=28.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W17 N$33 N$34 "Straight Waveguide" sch_x=1 sch_y=29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W18 N$35 N$36 "Straight Waveguide" sch_x=0 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W19 N$37 N$38 "Straight Waveguide" sch_x=4 sch_y=31.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W20 N$39 N$40 "Straight Waveguide" sch_x=3 sch_y=30.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W21 N$41 N$42 "Straight Waveguide" sch_x=3 sch_y=29.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W22 N$43 N$44 "Straight Waveguide" sch_x=5 sch_y=29.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W23 N$45 N$46 "Straight Waveguide" sch_x=5 sch_y=30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W24 N$47 N$48 "Straight Waveguide" sch_x=4 sch_y=28.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W25 N$49 N$50 "Straight Waveguide" sch_x=-4 sch_y=27.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W26 N$51 N$52 "Straight Waveguide" sch_x=-5 sch_y=26.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W27 N$53 N$54 "Straight Waveguide" sch_x=-5 sch_y=25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W28 N$55 N$56 "Straight Waveguide" sch_x=-3 sch_y=26.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W29 N$57 N$58 "Straight Waveguide" sch_x=-3 sch_y=25.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W30 N$59 N$60 "Straight Waveguide" sch_x=-4 sch_y=24.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W31 N$61 N$62 "Straight Waveguide" sch_x=0 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W32 N$63 N$64 "Straight Waveguide" sch_x=-1 sch_y=27.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W33 N$65 N$66 "Straight Waveguide" sch_x=-1 sch_y=26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W34 N$67 N$68 "Straight Waveguide" sch_x=1 sch_y=26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W35 N$69 N$70 "Straight Waveguide" sch_x=1 sch_y=27.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W36 N$71 N$72 "Straight Waveguide" sch_x=0 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W37 N$73 N$74 "Straight Waveguide" sch_x=0 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W38 N$75 N$76 "Straight Waveguide" sch_x=-1 sch_y=25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W39 N$77 N$78 "Straight Waveguide" sch_x=-1 sch_y=24.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W40 N$79 N$80 "Straight Waveguide" sch_x=1 sch_y=24.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W41 N$81 N$82 "Straight Waveguide" sch_x=1 sch_y=25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W42 N$83 N$84 "Straight Waveguide" sch_x=0 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W43 N$85 N$86 "Straight Waveguide" sch_x=4 sch_y=27.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W44 N$87 N$88 "Straight Waveguide" sch_x=3 sch_y=26.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W45 N$89 N$90 "Straight Waveguide" sch_x=3 sch_y=25.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W46 N$91 N$92 "Straight Waveguide" sch_x=5 sch_y=25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W47 N$93 N$94 "Straight Waveguide" sch_x=5 sch_y=26.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W48 N$95 N$96 "Straight Waveguide" sch_x=4 sch_y=24.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W49 N$98 N$97 "Straight Waveguide" sch_x=-13 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W50 N$100 N$99 "Straight Waveguide" sch_x=-13 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W51 N$102 N$101 "Straight Waveguide" sch_x=-13 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W52 N$104 N$103 "Straight Waveguide" sch_x=-13 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W53 N$106 N$105 "Straight Waveguide" sch_x=-13 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W54 N$108 N$107 "Straight Waveguide" sch_x=-13 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W55 N$110 N$109 "Straight Waveguide" sch_x=-11 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W56 N$112 N$111 "Straight Waveguide" sch_x=-11 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W57 N$114 N$113 "Straight Waveguide" sch_x=-11 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W58 N$116 N$115 "Straight Waveguide" sch_x=-11 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W59 N$118 N$117 "Straight Waveguide" sch_x=-9 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W60 N$120 N$119 "Straight Waveguide" sch_x=-9 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W61 N$121 N$122 "Straight Waveguide" sch_x=-9 sch_y=30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W62 N$123 N$124 "Straight Waveguide" sch_x=-8 sch_y=29.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W63 N$125 N$126 "Straight Waveguide" sch_x=-7 sch_y=28.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W64 N$127 N$128 "Straight Waveguide" sch_x=-7 sch_y=27.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W65 N$129 N$130 "Straight Waveguide" sch_x=-8 sch_y=26.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W66 N$131 N$132 "Straight Waveguide" sch_x=-9 sch_y=25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W67 N$133 N$134 "Straight Waveguide" sch_x=-10 sch_y=30.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W68 N$135 N$136 "Straight Waveguide" sch_x=-10 sch_y=25.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W69 N$137 N$138 "Straight Waveguide" sch_x=13 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W70 N$139 N$140 "Straight Waveguide" sch_x=13 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W71 N$141 N$142 "Straight Waveguide" sch_x=13 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W72 N$143 N$144 "Straight Waveguide" sch_x=13 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W73 N$145 N$146 "Straight Waveguide" sch_x=13 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W74 N$147 N$148 "Straight Waveguide" sch_x=13 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W75 N$149 N$150 "Straight Waveguide" sch_x=11 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W76 N$151 N$152 "Straight Waveguide" sch_x=11 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W77 N$153 N$154 "Straight Waveguide" sch_x=11 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W78 N$155 N$156 "Straight Waveguide" sch_x=11 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W79 N$157 N$158 "Straight Waveguide" sch_x=9 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W80 N$159 N$160 "Straight Waveguide" sch_x=9 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W81 N$162 N$161 "Straight Waveguide" sch_x=9 sch_y=30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W82 N$164 N$163 "Straight Waveguide" sch_x=8 sch_y=29.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W83 N$166 N$165 "Straight Waveguide" sch_x=7 sch_y=28.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W84 N$168 N$167 "Straight Waveguide" sch_x=7 sch_y=27.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W85 N$170 N$169 "Straight Waveguide" sch_x=8 sch_y=26.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W86 N$172 N$171 "Straight Waveguide" sch_x=9 sch_y=25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W87 N$174 N$173 "Straight Waveguide" sch_x=10 sch_y=30.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W88 N$176 N$175 "Straight Waveguide" sch_x=10 sch_y=25.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W89 N$177 N$178 "Straight Waveguide" sch_x=-4 sch_y=23.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W90 N$179 N$180 "Straight Waveguide" sch_x=-5 sch_y=22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W91 N$181 N$182 "Straight Waveguide" sch_x=-5 sch_y=21.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W92 N$183 N$184 "Straight Waveguide" sch_x=-3 sch_y=22.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W93 N$185 N$186 "Straight Waveguide" sch_x=-3 sch_y=21.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W94 N$187 N$188 "Straight Waveguide" sch_x=-4 sch_y=20.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W95 N$189 N$190 "Straight Waveguide" sch_x=0 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W96 N$191 N$192 "Straight Waveguide" sch_x=-1 sch_y=23.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W97 N$193 N$194 "Straight Waveguide" sch_x=-1 sch_y=22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W98 N$195 N$196 "Straight Waveguide" sch_x=1 sch_y=22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W99 N$197 N$198 "Straight Waveguide" sch_x=1 sch_y=23.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W100 N$199 N$200 "Straight Waveguide" sch_x=0 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W101 N$201 N$202 "Straight Waveguide" sch_x=0 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W102 N$203 N$204 "Straight Waveguide" sch_x=-1 sch_y=21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W103 N$205 N$206 "Straight Waveguide" sch_x=-1 sch_y=20.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W104 N$207 N$208 "Straight Waveguide" sch_x=1 sch_y=20.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W105 N$209 N$210 "Straight Waveguide" sch_x=1 sch_y=21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W106 N$211 N$212 "Straight Waveguide" sch_x=0 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W107 N$213 N$214 "Straight Waveguide" sch_x=4 sch_y=23.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W108 N$215 N$216 "Straight Waveguide" sch_x=3 sch_y=22.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W109 N$217 N$218 "Straight Waveguide" sch_x=3 sch_y=21.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W110 N$219 N$220 "Straight Waveguide" sch_x=5 sch_y=21.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W111 N$221 N$222 "Straight Waveguide" sch_x=5 sch_y=22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W112 N$223 N$224 "Straight Waveguide" sch_x=4 sch_y=20.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W113 N$225 N$226 "Straight Waveguide" sch_x=-4 sch_y=19.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W114 N$227 N$228 "Straight Waveguide" sch_x=-5 sch_y=18.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W115 N$229 N$230 "Straight Waveguide" sch_x=-5 sch_y=17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W116 N$231 N$232 "Straight Waveguide" sch_x=-3 sch_y=18.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W117 N$233 N$234 "Straight Waveguide" sch_x=-3 sch_y=17.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W118 N$235 N$236 "Straight Waveguide" sch_x=-4 sch_y=16.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W119 N$237 N$238 "Straight Waveguide" sch_x=0 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W120 N$239 N$240 "Straight Waveguide" sch_x=-1 sch_y=19.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W121 N$241 N$242 "Straight Waveguide" sch_x=-1 sch_y=18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W122 N$243 N$244 "Straight Waveguide" sch_x=1 sch_y=18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W123 N$245 N$246 "Straight Waveguide" sch_x=1 sch_y=19.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W124 N$247 N$248 "Straight Waveguide" sch_x=0 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W125 N$249 N$250 "Straight Waveguide" sch_x=0 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W126 N$251 N$252 "Straight Waveguide" sch_x=-1 sch_y=17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W127 N$253 N$254 "Straight Waveguide" sch_x=-1 sch_y=16.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W128 N$255 N$256 "Straight Waveguide" sch_x=1 sch_y=16.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W129 N$257 N$258 "Straight Waveguide" sch_x=1 sch_y=17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W130 N$259 N$260 "Straight Waveguide" sch_x=0 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W131 N$261 N$262 "Straight Waveguide" sch_x=4 sch_y=19.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W132 N$263 N$264 "Straight Waveguide" sch_x=3 sch_y=18.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W133 N$265 N$266 "Straight Waveguide" sch_x=3 sch_y=17.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W134 N$267 N$268 "Straight Waveguide" sch_x=5 sch_y=17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W135 N$269 N$270 "Straight Waveguide" sch_x=5 sch_y=18.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W136 N$271 N$272 "Straight Waveguide" sch_x=4 sch_y=16.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W137 N$274 N$273 "Straight Waveguide" sch_x=-13 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W138 N$276 N$275 "Straight Waveguide" sch_x=-13 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W139 N$278 N$277 "Straight Waveguide" sch_x=-13 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W140 N$280 N$279 "Straight Waveguide" sch_x=-13 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W141 N$282 N$281 "Straight Waveguide" sch_x=-13 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W142 N$284 N$283 "Straight Waveguide" sch_x=-13 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W143 N$286 N$285 "Straight Waveguide" sch_x=-11 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W144 N$288 N$287 "Straight Waveguide" sch_x=-11 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W145 N$290 N$289 "Straight Waveguide" sch_x=-11 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W146 N$292 N$291 "Straight Waveguide" sch_x=-11 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W147 N$294 N$293 "Straight Waveguide" sch_x=-9 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W148 N$296 N$295 "Straight Waveguide" sch_x=-9 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W149 N$297 N$298 "Straight Waveguide" sch_x=-9 sch_y=22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W150 N$299 N$300 "Straight Waveguide" sch_x=-8 sch_y=21.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W151 N$301 N$302 "Straight Waveguide" sch_x=-7 sch_y=20.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W152 N$303 N$304 "Straight Waveguide" sch_x=-7 sch_y=19.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W153 N$305 N$306 "Straight Waveguide" sch_x=-8 sch_y=18.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W154 N$307 N$308 "Straight Waveguide" sch_x=-9 sch_y=17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W155 N$309 N$310 "Straight Waveguide" sch_x=-10 sch_y=22.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W156 N$311 N$312 "Straight Waveguide" sch_x=-10 sch_y=17.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W157 N$313 N$314 "Straight Waveguide" sch_x=13 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W158 N$315 N$316 "Straight Waveguide" sch_x=13 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W159 N$317 N$318 "Straight Waveguide" sch_x=13 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W160 N$319 N$320 "Straight Waveguide" sch_x=13 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W161 N$321 N$322 "Straight Waveguide" sch_x=13 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W162 N$323 N$324 "Straight Waveguide" sch_x=13 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W163 N$325 N$326 "Straight Waveguide" sch_x=11 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W164 N$327 N$328 "Straight Waveguide" sch_x=11 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W165 N$329 N$330 "Straight Waveguide" sch_x=11 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W166 N$331 N$332 "Straight Waveguide" sch_x=11 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W167 N$333 N$334 "Straight Waveguide" sch_x=9 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W168 N$335 N$336 "Straight Waveguide" sch_x=9 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W169 N$338 N$337 "Straight Waveguide" sch_x=9 sch_y=22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W170 N$340 N$339 "Straight Waveguide" sch_x=8 sch_y=21.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W171 N$342 N$341 "Straight Waveguide" sch_x=7 sch_y=20.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W172 N$344 N$343 "Straight Waveguide" sch_x=7 sch_y=19.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W173 N$346 N$345 "Straight Waveguide" sch_x=8 sch_y=18.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W174 N$348 N$347 "Straight Waveguide" sch_x=9 sch_y=17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W175 N$350 N$349 "Straight Waveguide" sch_x=10 sch_y=22.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W176 N$352 N$351 "Straight Waveguide" sch_x=10 sch_y=17.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W177 N$354 N$353 "Straight Waveguide" sch_x=-29 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W178 N$356 N$355 "Straight Waveguide" sch_x=-29 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W179 N$358 N$357 "Straight Waveguide" sch_x=-29 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W180 N$360 N$359 "Straight Waveguide" sch_x=-29 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W181 N$362 N$361 "Straight Waveguide" sch_x=-29 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W182 N$364 N$363 "Straight Waveguide" sch_x=-29 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W183 N$366 N$365 "Straight Waveguide" sch_x=-29 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W184 N$368 N$367 "Straight Waveguide" sch_x=-29 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W185 N$370 N$369 "Straight Waveguide" sch_x=-29 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W186 N$372 N$371 "Straight Waveguide" sch_x=-29 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W187 N$374 N$373 "Straight Waveguide" sch_x=-29 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W188 N$376 N$375 "Straight Waveguide" sch_x=-29 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W189 N$378 N$377 "Straight Waveguide" sch_x=-29 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W190 N$380 N$379 "Straight Waveguide" sch_x=-29 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W191 N$382 N$381 "Straight Waveguide" sch_x=-27 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W192 N$384 N$383 "Straight Waveguide" sch_x=-27 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W193 N$386 N$385 "Straight Waveguide" sch_x=-27 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W194 N$388 N$387 "Straight Waveguide" sch_x=-27 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W195 N$390 N$389 "Straight Waveguide" sch_x=-27 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W196 N$392 N$391 "Straight Waveguide" sch_x=-27 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W197 N$394 N$393 "Straight Waveguide" sch_x=-27 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W198 N$396 N$395 "Straight Waveguide" sch_x=-27 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W199 N$398 N$397 "Straight Waveguide" sch_x=-27 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W200 N$400 N$399 "Straight Waveguide" sch_x=-27 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W201 N$402 N$401 "Straight Waveguide" sch_x=-27 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W202 N$404 N$403 "Straight Waveguide" sch_x=-27 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W203 N$406 N$405 "Straight Waveguide" sch_x=-25 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W204 N$408 N$407 "Straight Waveguide" sch_x=-25 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W205 N$410 N$409 "Straight Waveguide" sch_x=-25 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W206 N$412 N$411 "Straight Waveguide" sch_x=-25 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W207 N$414 N$413 "Straight Waveguide" sch_x=-25 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W208 N$416 N$415 "Straight Waveguide" sch_x=-25 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W209 N$418 N$417 "Straight Waveguide" sch_x=-25 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W210 N$420 N$419 "Straight Waveguide" sch_x=-25 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W211 N$422 N$421 "Straight Waveguide" sch_x=-25 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W212 N$424 N$423 "Straight Waveguide" sch_x=-25 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W213 N$426 N$425 "Straight Waveguide" sch_x=-23 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W214 N$428 N$427 "Straight Waveguide" sch_x=-23 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W215 N$430 N$429 "Straight Waveguide" sch_x=-23 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W216 N$432 N$431 "Straight Waveguide" sch_x=-23 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W217 N$434 N$433 "Straight Waveguide" sch_x=-23 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W218 N$436 N$435 "Straight Waveguide" sch_x=-23 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W219 N$438 N$437 "Straight Waveguide" sch_x=-23 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W220 N$440 N$439 "Straight Waveguide" sch_x=-23 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W221 N$442 N$441 "Straight Waveguide" sch_x=-21 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W222 N$444 N$443 "Straight Waveguide" sch_x=-21 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W223 N$446 N$445 "Straight Waveguide" sch_x=-21 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W224 N$448 N$447 "Straight Waveguide" sch_x=-21 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W225 N$450 N$449 "Straight Waveguide" sch_x=-21 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W226 N$452 N$451 "Straight Waveguide" sch_x=-21 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W227 N$454 N$453 "Straight Waveguide" sch_x=-19 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W228 N$456 N$455 "Straight Waveguide" sch_x=-19 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W229 N$458 N$457 "Straight Waveguide" sch_x=-19 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W230 N$460 N$459 "Straight Waveguide" sch_x=-19 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W231 N$462 N$461 "Straight Waveguide" sch_x=-17 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W232 N$464 N$463 "Straight Waveguide" sch_x=-17 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W233 N$465 N$466 "Straight Waveguide" sch_x=-21 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W234 N$467 N$468 "Straight Waveguide" sch_x=-20 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W235 N$469 N$470 "Straight Waveguide" sch_x=-19 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W236 N$471 N$472 "Straight Waveguide" sch_x=-18 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W237 N$473 N$474 "Straight Waveguide" sch_x=-17 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W238 N$475 N$476 "Straight Waveguide" sch_x=-16 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W239 N$477 N$478 "Straight Waveguide" sch_x=-15 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W240 N$479 N$480 "Straight Waveguide" sch_x=-15 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W241 N$481 N$482 "Straight Waveguide" sch_x=-16 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W242 N$483 N$484 "Straight Waveguide" sch_x=-17 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W243 N$485 N$486 "Straight Waveguide" sch_x=-18 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W244 N$487 N$488 "Straight Waveguide" sch_x=-19 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W245 N$489 N$490 "Straight Waveguide" sch_x=-20 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W246 N$491 N$492 "Straight Waveguide" sch_x=-21 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W247 N$493 N$494 "Straight Waveguide" sch_x=-22 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W248 N$495 N$496 "Straight Waveguide" sch_x=-22 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W249 N$497 N$498 "Straight Waveguide" sch_x=29 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W250 N$499 N$500 "Straight Waveguide" sch_x=29 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W251 N$501 N$502 "Straight Waveguide" sch_x=29 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W252 N$503 N$504 "Straight Waveguide" sch_x=29 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W253 N$505 N$506 "Straight Waveguide" sch_x=29 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W254 N$507 N$508 "Straight Waveguide" sch_x=29 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W255 N$509 N$510 "Straight Waveguide" sch_x=29 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W256 N$511 N$512 "Straight Waveguide" sch_x=29 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W257 N$513 N$514 "Straight Waveguide" sch_x=29 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W258 N$515 N$516 "Straight Waveguide" sch_x=29 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W259 N$517 N$518 "Straight Waveguide" sch_x=29 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W260 N$519 N$520 "Straight Waveguide" sch_x=29 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W261 N$521 N$522 "Straight Waveguide" sch_x=29 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W262 N$523 N$524 "Straight Waveguide" sch_x=29 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W263 N$525 N$526 "Straight Waveguide" sch_x=27 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W264 N$527 N$528 "Straight Waveguide" sch_x=27 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W265 N$529 N$530 "Straight Waveguide" sch_x=27 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W266 N$531 N$532 "Straight Waveguide" sch_x=27 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W267 N$533 N$534 "Straight Waveguide" sch_x=27 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W268 N$535 N$536 "Straight Waveguide" sch_x=27 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W269 N$537 N$538 "Straight Waveguide" sch_x=27 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W270 N$539 N$540 "Straight Waveguide" sch_x=27 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W271 N$541 N$542 "Straight Waveguide" sch_x=27 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W272 N$543 N$544 "Straight Waveguide" sch_x=27 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W273 N$545 N$546 "Straight Waveguide" sch_x=27 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W274 N$547 N$548 "Straight Waveguide" sch_x=27 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W275 N$549 N$550 "Straight Waveguide" sch_x=25 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W276 N$551 N$552 "Straight Waveguide" sch_x=25 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W277 N$553 N$554 "Straight Waveguide" sch_x=25 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W278 N$555 N$556 "Straight Waveguide" sch_x=25 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W279 N$557 N$558 "Straight Waveguide" sch_x=25 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W280 N$559 N$560 "Straight Waveguide" sch_x=25 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W281 N$561 N$562 "Straight Waveguide" sch_x=25 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W282 N$563 N$564 "Straight Waveguide" sch_x=25 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W283 N$565 N$566 "Straight Waveguide" sch_x=25 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W284 N$567 N$568 "Straight Waveguide" sch_x=25 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W285 N$569 N$570 "Straight Waveguide" sch_x=23 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W286 N$571 N$572 "Straight Waveguide" sch_x=23 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W287 N$573 N$574 "Straight Waveguide" sch_x=23 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W288 N$575 N$576 "Straight Waveguide" sch_x=23 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W289 N$577 N$578 "Straight Waveguide" sch_x=23 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W290 N$579 N$580 "Straight Waveguide" sch_x=23 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W291 N$581 N$582 "Straight Waveguide" sch_x=23 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W292 N$583 N$584 "Straight Waveguide" sch_x=23 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W293 N$585 N$586 "Straight Waveguide" sch_x=21 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W294 N$587 N$588 "Straight Waveguide" sch_x=21 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W295 N$589 N$590 "Straight Waveguide" sch_x=21 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W296 N$591 N$592 "Straight Waveguide" sch_x=21 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W297 N$593 N$594 "Straight Waveguide" sch_x=21 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W298 N$595 N$596 "Straight Waveguide" sch_x=21 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W299 N$597 N$598 "Straight Waveguide" sch_x=19 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W300 N$599 N$600 "Straight Waveguide" sch_x=19 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W301 N$601 N$602 "Straight Waveguide" sch_x=19 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W302 N$603 N$604 "Straight Waveguide" sch_x=19 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W303 N$605 N$606 "Straight Waveguide" sch_x=17 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W304 N$607 N$608 "Straight Waveguide" sch_x=17 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W305 N$610 N$609 "Straight Waveguide" sch_x=21 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W306 N$612 N$611 "Straight Waveguide" sch_x=20 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W307 N$614 N$613 "Straight Waveguide" sch_x=19 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W308 N$616 N$615 "Straight Waveguide" sch_x=18 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W309 N$618 N$617 "Straight Waveguide" sch_x=17 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W310 N$620 N$619 "Straight Waveguide" sch_x=16 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W311 N$622 N$621 "Straight Waveguide" sch_x=15 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W312 N$624 N$623 "Straight Waveguide" sch_x=15 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W313 N$626 N$625 "Straight Waveguide" sch_x=16 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W314 N$628 N$627 "Straight Waveguide" sch_x=17 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W315 N$630 N$629 "Straight Waveguide" sch_x=18 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W316 N$632 N$631 "Straight Waveguide" sch_x=19 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W317 N$634 N$633 "Straight Waveguide" sch_x=20 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W318 N$636 N$635 "Straight Waveguide" sch_x=21 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W319 N$638 N$637 "Straight Waveguide" sch_x=22 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W320 N$640 N$639 "Straight Waveguide" sch_x=22 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W321 N$641 N$642 "Straight Waveguide" sch_x=-4 sch_y=15.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W322 N$643 N$644 "Straight Waveguide" sch_x=-5 sch_y=14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W323 N$645 N$646 "Straight Waveguide" sch_x=-5 sch_y=13.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W324 N$647 N$648 "Straight Waveguide" sch_x=-3 sch_y=14.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W325 N$649 N$650 "Straight Waveguide" sch_x=-3 sch_y=13.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W326 N$651 N$652 "Straight Waveguide" sch_x=-4 sch_y=12.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W327 N$653 N$654 "Straight Waveguide" sch_x=0 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W328 N$655 N$656 "Straight Waveguide" sch_x=-1 sch_y=15.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W329 N$657 N$658 "Straight Waveguide" sch_x=-1 sch_y=14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W330 N$659 N$660 "Straight Waveguide" sch_x=1 sch_y=14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W331 N$661 N$662 "Straight Waveguide" sch_x=1 sch_y=15.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W332 N$663 N$664 "Straight Waveguide" sch_x=0 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W333 N$665 N$666 "Straight Waveguide" sch_x=0 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W334 N$667 N$668 "Straight Waveguide" sch_x=-1 sch_y=13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W335 N$669 N$670 "Straight Waveguide" sch_x=-1 sch_y=12.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W336 N$671 N$672 "Straight Waveguide" sch_x=1 sch_y=12.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W337 N$673 N$674 "Straight Waveguide" sch_x=1 sch_y=13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W338 N$675 N$676 "Straight Waveguide" sch_x=0 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W339 N$677 N$678 "Straight Waveguide" sch_x=4 sch_y=15.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W340 N$679 N$680 "Straight Waveguide" sch_x=3 sch_y=14.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W341 N$681 N$682 "Straight Waveguide" sch_x=3 sch_y=13.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W342 N$683 N$684 "Straight Waveguide" sch_x=5 sch_y=13.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W343 N$685 N$686 "Straight Waveguide" sch_x=5 sch_y=14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W344 N$687 N$688 "Straight Waveguide" sch_x=4 sch_y=12.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W345 N$689 N$690 "Straight Waveguide" sch_x=-4 sch_y=11.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W346 N$691 N$692 "Straight Waveguide" sch_x=-5 sch_y=10.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W347 N$693 N$694 "Straight Waveguide" sch_x=-5 sch_y=9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W348 N$695 N$696 "Straight Waveguide" sch_x=-3 sch_y=10.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W349 N$697 N$698 "Straight Waveguide" sch_x=-3 sch_y=9.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W350 N$699 N$700 "Straight Waveguide" sch_x=-4 sch_y=8.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W351 N$701 N$702 "Straight Waveguide" sch_x=0 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W352 N$703 N$704 "Straight Waveguide" sch_x=-1 sch_y=11.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W353 N$705 N$706 "Straight Waveguide" sch_x=-1 sch_y=10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W354 N$707 N$708 "Straight Waveguide" sch_x=1 sch_y=10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W355 N$709 N$710 "Straight Waveguide" sch_x=1 sch_y=11.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W356 N$711 N$712 "Straight Waveguide" sch_x=0 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W357 N$713 N$714 "Straight Waveguide" sch_x=0 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W358 N$715 N$716 "Straight Waveguide" sch_x=-1 sch_y=9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W359 N$717 N$718 "Straight Waveguide" sch_x=-1 sch_y=8.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W360 N$719 N$720 "Straight Waveguide" sch_x=1 sch_y=8.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W361 N$721 N$722 "Straight Waveguide" sch_x=1 sch_y=9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W362 N$723 N$724 "Straight Waveguide" sch_x=0 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W363 N$725 N$726 "Straight Waveguide" sch_x=4 sch_y=11.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W364 N$727 N$728 "Straight Waveguide" sch_x=3 sch_y=10.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W365 N$729 N$730 "Straight Waveguide" sch_x=3 sch_y=9.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W366 N$731 N$732 "Straight Waveguide" sch_x=5 sch_y=9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W367 N$733 N$734 "Straight Waveguide" sch_x=5 sch_y=10.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W368 N$735 N$736 "Straight Waveguide" sch_x=4 sch_y=8.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W369 N$738 N$737 "Straight Waveguide" sch_x=-13 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W370 N$740 N$739 "Straight Waveguide" sch_x=-13 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W371 N$742 N$741 "Straight Waveguide" sch_x=-13 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W372 N$744 N$743 "Straight Waveguide" sch_x=-13 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W373 N$746 N$745 "Straight Waveguide" sch_x=-13 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W374 N$748 N$747 "Straight Waveguide" sch_x=-13 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W375 N$750 N$749 "Straight Waveguide" sch_x=-11 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W376 N$752 N$751 "Straight Waveguide" sch_x=-11 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W377 N$754 N$753 "Straight Waveguide" sch_x=-11 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W378 N$756 N$755 "Straight Waveguide" sch_x=-11 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W379 N$758 N$757 "Straight Waveguide" sch_x=-9 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W380 N$760 N$759 "Straight Waveguide" sch_x=-9 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W381 N$761 N$762 "Straight Waveguide" sch_x=-9 sch_y=14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W382 N$763 N$764 "Straight Waveguide" sch_x=-8 sch_y=13.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W383 N$765 N$766 "Straight Waveguide" sch_x=-7 sch_y=12.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W384 N$767 N$768 "Straight Waveguide" sch_x=-7 sch_y=11.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W385 N$769 N$770 "Straight Waveguide" sch_x=-8 sch_y=10.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W386 N$771 N$772 "Straight Waveguide" sch_x=-9 sch_y=9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W387 N$773 N$774 "Straight Waveguide" sch_x=-10 sch_y=14.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W388 N$775 N$776 "Straight Waveguide" sch_x=-10 sch_y=9.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W389 N$777 N$778 "Straight Waveguide" sch_x=13 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W390 N$779 N$780 "Straight Waveguide" sch_x=13 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W391 N$781 N$782 "Straight Waveguide" sch_x=13 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W392 N$783 N$784 "Straight Waveguide" sch_x=13 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W393 N$785 N$786 "Straight Waveguide" sch_x=13 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W394 N$787 N$788 "Straight Waveguide" sch_x=13 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W395 N$789 N$790 "Straight Waveguide" sch_x=11 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W396 N$791 N$792 "Straight Waveguide" sch_x=11 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W397 N$793 N$794 "Straight Waveguide" sch_x=11 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W398 N$795 N$796 "Straight Waveguide" sch_x=11 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W399 N$797 N$798 "Straight Waveguide" sch_x=9 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W400 N$799 N$800 "Straight Waveguide" sch_x=9 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W401 N$802 N$801 "Straight Waveguide" sch_x=9 sch_y=14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W402 N$804 N$803 "Straight Waveguide" sch_x=8 sch_y=13.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W403 N$806 N$805 "Straight Waveguide" sch_x=7 sch_y=12.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W404 N$808 N$807 "Straight Waveguide" sch_x=7 sch_y=11.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W405 N$810 N$809 "Straight Waveguide" sch_x=8 sch_y=10.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W406 N$812 N$811 "Straight Waveguide" sch_x=9 sch_y=9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W407 N$814 N$813 "Straight Waveguide" sch_x=10 sch_y=14.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W408 N$816 N$815 "Straight Waveguide" sch_x=10 sch_y=9.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W409 N$817 N$818 "Straight Waveguide" sch_x=-4 sch_y=7.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W410 N$819 N$820 "Straight Waveguide" sch_x=-5 sch_y=6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W411 N$821 N$822 "Straight Waveguide" sch_x=-5 sch_y=5.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W412 N$823 N$824 "Straight Waveguide" sch_x=-3 sch_y=6.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W413 N$825 N$826 "Straight Waveguide" sch_x=-3 sch_y=5.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W414 N$827 N$828 "Straight Waveguide" sch_x=-4 sch_y=4.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W415 N$829 N$830 "Straight Waveguide" sch_x=0 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W416 N$831 N$832 "Straight Waveguide" sch_x=-1 sch_y=7.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W417 N$833 N$834 "Straight Waveguide" sch_x=-1 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W418 N$835 N$836 "Straight Waveguide" sch_x=1 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W419 N$837 N$838 "Straight Waveguide" sch_x=1 sch_y=7.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W420 N$839 N$840 "Straight Waveguide" sch_x=0 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W421 N$841 N$842 "Straight Waveguide" sch_x=0 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W422 N$843 N$844 "Straight Waveguide" sch_x=-1 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W423 N$845 N$846 "Straight Waveguide" sch_x=-1 sch_y=4.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W424 N$847 N$848 "Straight Waveguide" sch_x=1 sch_y=4.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W425 N$849 N$850 "Straight Waveguide" sch_x=1 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W426 N$851 N$852 "Straight Waveguide" sch_x=0 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W427 N$853 N$854 "Straight Waveguide" sch_x=4 sch_y=7.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W428 N$855 N$856 "Straight Waveguide" sch_x=3 sch_y=6.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W429 N$857 N$858 "Straight Waveguide" sch_x=3 sch_y=5.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W430 N$859 N$860 "Straight Waveguide" sch_x=5 sch_y=5.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W431 N$861 N$862 "Straight Waveguide" sch_x=5 sch_y=6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W432 N$863 N$864 "Straight Waveguide" sch_x=4 sch_y=4.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W433 N$865 N$866 "Straight Waveguide" sch_x=-4 sch_y=3.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W434 N$867 N$868 "Straight Waveguide" sch_x=-5 sch_y=2.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W435 N$869 N$870 "Straight Waveguide" sch_x=-5 sch_y=1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W436 N$871 N$872 "Straight Waveguide" sch_x=-3 sch_y=2.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W437 N$873 N$874 "Straight Waveguide" sch_x=-3 sch_y=1.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W438 N$875 N$876 "Straight Waveguide" sch_x=-4 sch_y=0.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W439 N$877 N$878 "Straight Waveguide" sch_x=0 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W440 N$879 N$880 "Straight Waveguide" sch_x=-1 sch_y=3.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W441 N$881 N$882 "Straight Waveguide" sch_x=-1 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W442 N$883 N$884 "Straight Waveguide" sch_x=1 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W443 N$885 N$886 "Straight Waveguide" sch_x=1 sch_y=3.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W444 N$887 N$888 "Straight Waveguide" sch_x=0 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W445 N$889 N$890 "Straight Waveguide" sch_x=0 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W446 N$891 N$892 "Straight Waveguide" sch_x=-1 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W447 N$893 N$894 "Straight Waveguide" sch_x=-1 sch_y=0.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W448 N$895 N$896 "Straight Waveguide" sch_x=1 sch_y=0.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W449 N$897 N$898 "Straight Waveguide" sch_x=1 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W450 N$899 N$900 "Straight Waveguide" sch_x=0 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W451 N$901 N$902 "Straight Waveguide" sch_x=4 sch_y=3.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W452 N$903 N$904 "Straight Waveguide" sch_x=3 sch_y=2.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W453 N$905 N$906 "Straight Waveguide" sch_x=3 sch_y=1.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W454 N$907 N$908 "Straight Waveguide" sch_x=5 sch_y=1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W455 N$909 N$910 "Straight Waveguide" sch_x=5 sch_y=2.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W456 N$911 N$912 "Straight Waveguide" sch_x=4 sch_y=0.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W457 N$914 N$913 "Straight Waveguide" sch_x=-13 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W458 N$916 N$915 "Straight Waveguide" sch_x=-13 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W459 N$918 N$917 "Straight Waveguide" sch_x=-13 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W460 N$920 N$919 "Straight Waveguide" sch_x=-13 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W461 N$922 N$921 "Straight Waveguide" sch_x=-13 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W462 N$924 N$923 "Straight Waveguide" sch_x=-13 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W463 N$926 N$925 "Straight Waveguide" sch_x=-11 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W464 N$928 N$927 "Straight Waveguide" sch_x=-11 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W465 N$930 N$929 "Straight Waveguide" sch_x=-11 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W466 N$932 N$931 "Straight Waveguide" sch_x=-11 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W467 N$934 N$933 "Straight Waveguide" sch_x=-9 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W468 N$936 N$935 "Straight Waveguide" sch_x=-9 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W469 N$937 N$938 "Straight Waveguide" sch_x=-9 sch_y=6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W470 N$939 N$940 "Straight Waveguide" sch_x=-8 sch_y=5.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W471 N$941 N$942 "Straight Waveguide" sch_x=-7 sch_y=4.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W472 N$943 N$944 "Straight Waveguide" sch_x=-7 sch_y=3.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W473 N$945 N$946 "Straight Waveguide" sch_x=-8 sch_y=2.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W474 N$947 N$948 "Straight Waveguide" sch_x=-9 sch_y=1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W475 N$949 N$950 "Straight Waveguide" sch_x=-10 sch_y=6.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W476 N$951 N$952 "Straight Waveguide" sch_x=-10 sch_y=1.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W477 N$953 N$954 "Straight Waveguide" sch_x=13 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W478 N$955 N$956 "Straight Waveguide" sch_x=13 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W479 N$957 N$958 "Straight Waveguide" sch_x=13 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W480 N$959 N$960 "Straight Waveguide" sch_x=13 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W481 N$961 N$962 "Straight Waveguide" sch_x=13 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W482 N$963 N$964 "Straight Waveguide" sch_x=13 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W483 N$965 N$966 "Straight Waveguide" sch_x=11 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W484 N$967 N$968 "Straight Waveguide" sch_x=11 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W485 N$969 N$970 "Straight Waveguide" sch_x=11 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W486 N$971 N$972 "Straight Waveguide" sch_x=11 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W487 N$973 N$974 "Straight Waveguide" sch_x=9 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W488 N$975 N$976 "Straight Waveguide" sch_x=9 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W489 N$978 N$977 "Straight Waveguide" sch_x=9 sch_y=6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W490 N$980 N$979 "Straight Waveguide" sch_x=8 sch_y=5.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W491 N$982 N$981 "Straight Waveguide" sch_x=7 sch_y=4.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W492 N$984 N$983 "Straight Waveguide" sch_x=7 sch_y=3.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W493 N$986 N$985 "Straight Waveguide" sch_x=8 sch_y=2.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W494 N$988 N$987 "Straight Waveguide" sch_x=9 sch_y=1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W495 N$990 N$989 "Straight Waveguide" sch_x=10 sch_y=6.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W496 N$992 N$991 "Straight Waveguide" sch_x=10 sch_y=1.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W497 N$994 N$993 "Straight Waveguide" sch_x=-29 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W498 N$996 N$995 "Straight Waveguide" sch_x=-29 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W499 N$998 N$997 "Straight Waveguide" sch_x=-29 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W500 N$1000 N$999 "Straight Waveguide" sch_x=-29 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W501 N$1002 N$1001 "Straight Waveguide" sch_x=-29 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W502 N$1004 N$1003 "Straight Waveguide" sch_x=-29 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W503 N$1006 N$1005 "Straight Waveguide" sch_x=-29 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W504 N$1008 N$1007 "Straight Waveguide" sch_x=-29 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W505 N$1010 N$1009 "Straight Waveguide" sch_x=-29 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W506 N$1012 N$1011 "Straight Waveguide" sch_x=-29 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W507 N$1014 N$1013 "Straight Waveguide" sch_x=-29 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W508 N$1016 N$1015 "Straight Waveguide" sch_x=-29 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W509 N$1018 N$1017 "Straight Waveguide" sch_x=-29 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W510 N$1020 N$1019 "Straight Waveguide" sch_x=-29 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W511 N$1022 N$1021 "Straight Waveguide" sch_x=-27 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W512 N$1024 N$1023 "Straight Waveguide" sch_x=-27 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W513 N$1026 N$1025 "Straight Waveguide" sch_x=-27 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W514 N$1028 N$1027 "Straight Waveguide" sch_x=-27 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W515 N$1030 N$1029 "Straight Waveguide" sch_x=-27 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W516 N$1032 N$1031 "Straight Waveguide" sch_x=-27 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W517 N$1034 N$1033 "Straight Waveguide" sch_x=-27 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W518 N$1036 N$1035 "Straight Waveguide" sch_x=-27 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W519 N$1038 N$1037 "Straight Waveguide" sch_x=-27 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W520 N$1040 N$1039 "Straight Waveguide" sch_x=-27 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W521 N$1042 N$1041 "Straight Waveguide" sch_x=-27 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W522 N$1044 N$1043 "Straight Waveguide" sch_x=-27 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W523 N$1046 N$1045 "Straight Waveguide" sch_x=-25 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W524 N$1048 N$1047 "Straight Waveguide" sch_x=-25 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W525 N$1050 N$1049 "Straight Waveguide" sch_x=-25 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W526 N$1052 N$1051 "Straight Waveguide" sch_x=-25 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W527 N$1054 N$1053 "Straight Waveguide" sch_x=-25 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W528 N$1056 N$1055 "Straight Waveguide" sch_x=-25 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W529 N$1058 N$1057 "Straight Waveguide" sch_x=-25 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W530 N$1060 N$1059 "Straight Waveguide" sch_x=-25 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W531 N$1062 N$1061 "Straight Waveguide" sch_x=-25 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W532 N$1064 N$1063 "Straight Waveguide" sch_x=-25 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W533 N$1066 N$1065 "Straight Waveguide" sch_x=-23 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W534 N$1068 N$1067 "Straight Waveguide" sch_x=-23 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W535 N$1070 N$1069 "Straight Waveguide" sch_x=-23 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W536 N$1072 N$1071 "Straight Waveguide" sch_x=-23 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W537 N$1074 N$1073 "Straight Waveguide" sch_x=-23 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W538 N$1076 N$1075 "Straight Waveguide" sch_x=-23 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W539 N$1078 N$1077 "Straight Waveguide" sch_x=-23 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W540 N$1080 N$1079 "Straight Waveguide" sch_x=-23 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W541 N$1082 N$1081 "Straight Waveguide" sch_x=-21 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W542 N$1084 N$1083 "Straight Waveguide" sch_x=-21 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W543 N$1086 N$1085 "Straight Waveguide" sch_x=-21 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W544 N$1088 N$1087 "Straight Waveguide" sch_x=-21 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W545 N$1090 N$1089 "Straight Waveguide" sch_x=-21 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W546 N$1092 N$1091 "Straight Waveguide" sch_x=-21 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W547 N$1094 N$1093 "Straight Waveguide" sch_x=-19 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W548 N$1096 N$1095 "Straight Waveguide" sch_x=-19 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W549 N$1098 N$1097 "Straight Waveguide" sch_x=-19 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W550 N$1100 N$1099 "Straight Waveguide" sch_x=-19 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W551 N$1102 N$1101 "Straight Waveguide" sch_x=-17 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W552 N$1104 N$1103 "Straight Waveguide" sch_x=-17 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W553 N$1105 N$1106 "Straight Waveguide" sch_x=-21 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W554 N$1107 N$1108 "Straight Waveguide" sch_x=-20 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W555 N$1109 N$1110 "Straight Waveguide" sch_x=-19 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W556 N$1111 N$1112 "Straight Waveguide" sch_x=-18 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W557 N$1113 N$1114 "Straight Waveguide" sch_x=-17 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W558 N$1115 N$1116 "Straight Waveguide" sch_x=-16 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W559 N$1117 N$1118 "Straight Waveguide" sch_x=-15 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W560 N$1119 N$1120 "Straight Waveguide" sch_x=-15 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W561 N$1121 N$1122 "Straight Waveguide" sch_x=-16 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W562 N$1123 N$1124 "Straight Waveguide" sch_x=-17 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W563 N$1125 N$1126 "Straight Waveguide" sch_x=-18 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W564 N$1127 N$1128 "Straight Waveguide" sch_x=-19 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W565 N$1129 N$1130 "Straight Waveguide" sch_x=-20 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W566 N$1131 N$1132 "Straight Waveguide" sch_x=-21 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W567 N$1133 N$1134 "Straight Waveguide" sch_x=-22 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W568 N$1135 N$1136 "Straight Waveguide" sch_x=-22 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W569 N$1137 N$1138 "Straight Waveguide" sch_x=29 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W570 N$1139 N$1140 "Straight Waveguide" sch_x=29 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W571 N$1141 N$1142 "Straight Waveguide" sch_x=29 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W572 N$1143 N$1144 "Straight Waveguide" sch_x=29 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W573 N$1145 N$1146 "Straight Waveguide" sch_x=29 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W574 N$1147 N$1148 "Straight Waveguide" sch_x=29 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W575 N$1149 N$1150 "Straight Waveguide" sch_x=29 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W576 N$1151 N$1152 "Straight Waveguide" sch_x=29 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W577 N$1153 N$1154 "Straight Waveguide" sch_x=29 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W578 N$1155 N$1156 "Straight Waveguide" sch_x=29 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W579 N$1157 N$1158 "Straight Waveguide" sch_x=29 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W580 N$1159 N$1160 "Straight Waveguide" sch_x=29 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W581 N$1161 N$1162 "Straight Waveguide" sch_x=29 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W582 N$1163 N$1164 "Straight Waveguide" sch_x=29 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W583 N$1165 N$1166 "Straight Waveguide" sch_x=27 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W584 N$1167 N$1168 "Straight Waveguide" sch_x=27 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W585 N$1169 N$1170 "Straight Waveguide" sch_x=27 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W586 N$1171 N$1172 "Straight Waveguide" sch_x=27 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W587 N$1173 N$1174 "Straight Waveguide" sch_x=27 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W588 N$1175 N$1176 "Straight Waveguide" sch_x=27 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W589 N$1177 N$1178 "Straight Waveguide" sch_x=27 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W590 N$1179 N$1180 "Straight Waveguide" sch_x=27 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W591 N$1181 N$1182 "Straight Waveguide" sch_x=27 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W592 N$1183 N$1184 "Straight Waveguide" sch_x=27 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W593 N$1185 N$1186 "Straight Waveguide" sch_x=27 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W594 N$1187 N$1188 "Straight Waveguide" sch_x=27 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W595 N$1189 N$1190 "Straight Waveguide" sch_x=25 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W596 N$1191 N$1192 "Straight Waveguide" sch_x=25 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W597 N$1193 N$1194 "Straight Waveguide" sch_x=25 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W598 N$1195 N$1196 "Straight Waveguide" sch_x=25 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W599 N$1197 N$1198 "Straight Waveguide" sch_x=25 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W600 N$1199 N$1200 "Straight Waveguide" sch_x=25 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W601 N$1201 N$1202 "Straight Waveguide" sch_x=25 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W602 N$1203 N$1204 "Straight Waveguide" sch_x=25 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W603 N$1205 N$1206 "Straight Waveguide" sch_x=25 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W604 N$1207 N$1208 "Straight Waveguide" sch_x=25 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W605 N$1209 N$1210 "Straight Waveguide" sch_x=23 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W606 N$1211 N$1212 "Straight Waveguide" sch_x=23 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W607 N$1213 N$1214 "Straight Waveguide" sch_x=23 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W608 N$1215 N$1216 "Straight Waveguide" sch_x=23 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W609 N$1217 N$1218 "Straight Waveguide" sch_x=23 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W610 N$1219 N$1220 "Straight Waveguide" sch_x=23 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W611 N$1221 N$1222 "Straight Waveguide" sch_x=23 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W612 N$1223 N$1224 "Straight Waveguide" sch_x=23 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W613 N$1225 N$1226 "Straight Waveguide" sch_x=21 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W614 N$1227 N$1228 "Straight Waveguide" sch_x=21 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W615 N$1229 N$1230 "Straight Waveguide" sch_x=21 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W616 N$1231 N$1232 "Straight Waveguide" sch_x=21 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W617 N$1233 N$1234 "Straight Waveguide" sch_x=21 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W618 N$1235 N$1236 "Straight Waveguide" sch_x=21 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W619 N$1237 N$1238 "Straight Waveguide" sch_x=19 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W620 N$1239 N$1240 "Straight Waveguide" sch_x=19 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W621 N$1241 N$1242 "Straight Waveguide" sch_x=19 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W622 N$1243 N$1244 "Straight Waveguide" sch_x=19 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W623 N$1245 N$1246 "Straight Waveguide" sch_x=17 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W624 N$1247 N$1248 "Straight Waveguide" sch_x=17 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W625 N$1250 N$1249 "Straight Waveguide" sch_x=21 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W626 N$1252 N$1251 "Straight Waveguide" sch_x=20 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W627 N$1254 N$1253 "Straight Waveguide" sch_x=19 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W628 N$1256 N$1255 "Straight Waveguide" sch_x=18 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W629 N$1258 N$1257 "Straight Waveguide" sch_x=17 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W630 N$1260 N$1259 "Straight Waveguide" sch_x=16 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W631 N$1262 N$1261 "Straight Waveguide" sch_x=15 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W632 N$1264 N$1263 "Straight Waveguide" sch_x=15 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W633 N$1266 N$1265 "Straight Waveguide" sch_x=16 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W634 N$1268 N$1267 "Straight Waveguide" sch_x=17 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W635 N$1270 N$1269 "Straight Waveguide" sch_x=18 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W636 N$1272 N$1271 "Straight Waveguide" sch_x=19 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W637 N$1274 N$1273 "Straight Waveguide" sch_x=20 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W638 N$1276 N$1275 "Straight Waveguide" sch_x=21 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W639 N$1278 N$1277 "Straight Waveguide" sch_x=22 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W640 N$1280 N$1279 "Straight Waveguide" sch_x=22 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W641 N$1282 N$1281 "Straight Waveguide" sch_x=-61 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W642 N$1284 N$1283 "Straight Waveguide" sch_x=-61 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W643 N$1286 N$1285 "Straight Waveguide" sch_x=-61 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W644 N$1288 N$1287 "Straight Waveguide" sch_x=-61 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W645 N$1290 N$1289 "Straight Waveguide" sch_x=-61 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W646 N$1292 N$1291 "Straight Waveguide" sch_x=-61 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W647 N$1294 N$1293 "Straight Waveguide" sch_x=-61 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W648 N$1296 N$1295 "Straight Waveguide" sch_x=-61 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W649 N$1298 N$1297 "Straight Waveguide" sch_x=-61 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W650 N$1300 N$1299 "Straight Waveguide" sch_x=-61 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W651 N$1302 N$1301 "Straight Waveguide" sch_x=-61 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W652 N$1304 N$1303 "Straight Waveguide" sch_x=-61 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W653 N$1306 N$1305 "Straight Waveguide" sch_x=-61 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W654 N$1308 N$1307 "Straight Waveguide" sch_x=-61 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W655 N$1310 N$1309 "Straight Waveguide" sch_x=-61 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W656 N$1312 N$1311 "Straight Waveguide" sch_x=-61 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W657 N$1314 N$1313 "Straight Waveguide" sch_x=-61 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W658 N$1316 N$1315 "Straight Waveguide" sch_x=-61 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W659 N$1318 N$1317 "Straight Waveguide" sch_x=-61 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W660 N$1320 N$1319 "Straight Waveguide" sch_x=-61 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W661 N$1322 N$1321 "Straight Waveguide" sch_x=-61 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W662 N$1324 N$1323 "Straight Waveguide" sch_x=-61 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W663 N$1326 N$1325 "Straight Waveguide" sch_x=-61 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W664 N$1328 N$1327 "Straight Waveguide" sch_x=-61 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W665 N$1330 N$1329 "Straight Waveguide" sch_x=-61 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W666 N$1332 N$1331 "Straight Waveguide" sch_x=-61 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W667 N$1334 N$1333 "Straight Waveguide" sch_x=-61 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W668 N$1336 N$1335 "Straight Waveguide" sch_x=-61 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W669 N$1338 N$1337 "Straight Waveguide" sch_x=-61 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W670 N$1340 N$1339 "Straight Waveguide" sch_x=-61 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W671 N$1342 N$1341 "Straight Waveguide" sch_x=-59 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W672 N$1344 N$1343 "Straight Waveguide" sch_x=-59 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W673 N$1346 N$1345 "Straight Waveguide" sch_x=-59 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W674 N$1348 N$1347 "Straight Waveguide" sch_x=-59 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W675 N$1350 N$1349 "Straight Waveguide" sch_x=-59 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W676 N$1352 N$1351 "Straight Waveguide" sch_x=-59 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W677 N$1354 N$1353 "Straight Waveguide" sch_x=-59 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W678 N$1356 N$1355 "Straight Waveguide" sch_x=-59 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W679 N$1358 N$1357 "Straight Waveguide" sch_x=-59 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W680 N$1360 N$1359 "Straight Waveguide" sch_x=-59 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W681 N$1362 N$1361 "Straight Waveguide" sch_x=-59 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W682 N$1364 N$1363 "Straight Waveguide" sch_x=-59 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W683 N$1366 N$1365 "Straight Waveguide" sch_x=-59 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W684 N$1368 N$1367 "Straight Waveguide" sch_x=-59 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W685 N$1370 N$1369 "Straight Waveguide" sch_x=-59 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W686 N$1372 N$1371 "Straight Waveguide" sch_x=-59 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W687 N$1374 N$1373 "Straight Waveguide" sch_x=-59 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W688 N$1376 N$1375 "Straight Waveguide" sch_x=-59 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W689 N$1378 N$1377 "Straight Waveguide" sch_x=-59 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W690 N$1380 N$1379 "Straight Waveguide" sch_x=-59 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W691 N$1382 N$1381 "Straight Waveguide" sch_x=-59 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W692 N$1384 N$1383 "Straight Waveguide" sch_x=-59 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W693 N$1386 N$1385 "Straight Waveguide" sch_x=-59 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W694 N$1388 N$1387 "Straight Waveguide" sch_x=-59 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W695 N$1390 N$1389 "Straight Waveguide" sch_x=-59 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W696 N$1392 N$1391 "Straight Waveguide" sch_x=-59 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W697 N$1394 N$1393 "Straight Waveguide" sch_x=-59 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W698 N$1396 N$1395 "Straight Waveguide" sch_x=-59 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W699 N$1398 N$1397 "Straight Waveguide" sch_x=-57 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W700 N$1400 N$1399 "Straight Waveguide" sch_x=-57 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W701 N$1402 N$1401 "Straight Waveguide" sch_x=-57 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W702 N$1404 N$1403 "Straight Waveguide" sch_x=-57 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W703 N$1406 N$1405 "Straight Waveguide" sch_x=-57 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W704 N$1408 N$1407 "Straight Waveguide" sch_x=-57 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W705 N$1410 N$1409 "Straight Waveguide" sch_x=-57 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W706 N$1412 N$1411 "Straight Waveguide" sch_x=-57 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W707 N$1414 N$1413 "Straight Waveguide" sch_x=-57 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W708 N$1416 N$1415 "Straight Waveguide" sch_x=-57 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W709 N$1418 N$1417 "Straight Waveguide" sch_x=-57 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W710 N$1420 N$1419 "Straight Waveguide" sch_x=-57 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W711 N$1422 N$1421 "Straight Waveguide" sch_x=-57 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W712 N$1424 N$1423 "Straight Waveguide" sch_x=-57 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W713 N$1426 N$1425 "Straight Waveguide" sch_x=-57 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W714 N$1428 N$1427 "Straight Waveguide" sch_x=-57 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W715 N$1430 N$1429 "Straight Waveguide" sch_x=-57 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W716 N$1432 N$1431 "Straight Waveguide" sch_x=-57 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W717 N$1434 N$1433 "Straight Waveguide" sch_x=-57 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W718 N$1436 N$1435 "Straight Waveguide" sch_x=-57 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W719 N$1438 N$1437 "Straight Waveguide" sch_x=-57 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W720 N$1440 N$1439 "Straight Waveguide" sch_x=-57 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W721 N$1442 N$1441 "Straight Waveguide" sch_x=-57 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W722 N$1444 N$1443 "Straight Waveguide" sch_x=-57 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W723 N$1446 N$1445 "Straight Waveguide" sch_x=-57 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W724 N$1448 N$1447 "Straight Waveguide" sch_x=-57 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W725 N$1450 N$1449 "Straight Waveguide" sch_x=-55 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W726 N$1452 N$1451 "Straight Waveguide" sch_x=-55 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W727 N$1454 N$1453 "Straight Waveguide" sch_x=-55 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W728 N$1456 N$1455 "Straight Waveguide" sch_x=-55 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W729 N$1458 N$1457 "Straight Waveguide" sch_x=-55 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W730 N$1460 N$1459 "Straight Waveguide" sch_x=-55 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W731 N$1462 N$1461 "Straight Waveguide" sch_x=-55 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W732 N$1464 N$1463 "Straight Waveguide" sch_x=-55 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W733 N$1466 N$1465 "Straight Waveguide" sch_x=-55 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W734 N$1468 N$1467 "Straight Waveguide" sch_x=-55 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W735 N$1470 N$1469 "Straight Waveguide" sch_x=-55 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W736 N$1472 N$1471 "Straight Waveguide" sch_x=-55 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W737 N$1474 N$1473 "Straight Waveguide" sch_x=-55 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W738 N$1476 N$1475 "Straight Waveguide" sch_x=-55 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W739 N$1478 N$1477 "Straight Waveguide" sch_x=-55 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W740 N$1480 N$1479 "Straight Waveguide" sch_x=-55 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W741 N$1482 N$1481 "Straight Waveguide" sch_x=-55 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W742 N$1484 N$1483 "Straight Waveguide" sch_x=-55 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W743 N$1486 N$1485 "Straight Waveguide" sch_x=-55 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W744 N$1488 N$1487 "Straight Waveguide" sch_x=-55 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W745 N$1490 N$1489 "Straight Waveguide" sch_x=-55 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W746 N$1492 N$1491 "Straight Waveguide" sch_x=-55 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W747 N$1494 N$1493 "Straight Waveguide" sch_x=-55 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W748 N$1496 N$1495 "Straight Waveguide" sch_x=-55 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W749 N$1498 N$1497 "Straight Waveguide" sch_x=-53 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W750 N$1500 N$1499 "Straight Waveguide" sch_x=-53 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W751 N$1502 N$1501 "Straight Waveguide" sch_x=-53 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W752 N$1504 N$1503 "Straight Waveguide" sch_x=-53 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W753 N$1506 N$1505 "Straight Waveguide" sch_x=-53 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W754 N$1508 N$1507 "Straight Waveguide" sch_x=-53 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W755 N$1510 N$1509 "Straight Waveguide" sch_x=-53 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W756 N$1512 N$1511 "Straight Waveguide" sch_x=-53 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W757 N$1514 N$1513 "Straight Waveguide" sch_x=-53 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W758 N$1516 N$1515 "Straight Waveguide" sch_x=-53 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W759 N$1518 N$1517 "Straight Waveguide" sch_x=-53 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W760 N$1520 N$1519 "Straight Waveguide" sch_x=-53 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W761 N$1522 N$1521 "Straight Waveguide" sch_x=-53 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W762 N$1524 N$1523 "Straight Waveguide" sch_x=-53 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W763 N$1526 N$1525 "Straight Waveguide" sch_x=-53 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W764 N$1528 N$1527 "Straight Waveguide" sch_x=-53 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W765 N$1530 N$1529 "Straight Waveguide" sch_x=-53 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W766 N$1532 N$1531 "Straight Waveguide" sch_x=-53 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W767 N$1534 N$1533 "Straight Waveguide" sch_x=-53 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W768 N$1536 N$1535 "Straight Waveguide" sch_x=-53 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W769 N$1538 N$1537 "Straight Waveguide" sch_x=-53 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W770 N$1540 N$1539 "Straight Waveguide" sch_x=-53 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W771 N$1542 N$1541 "Straight Waveguide" sch_x=-51 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W772 N$1544 N$1543 "Straight Waveguide" sch_x=-51 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W773 N$1546 N$1545 "Straight Waveguide" sch_x=-51 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W774 N$1548 N$1547 "Straight Waveguide" sch_x=-51 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W775 N$1550 N$1549 "Straight Waveguide" sch_x=-51 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W776 N$1552 N$1551 "Straight Waveguide" sch_x=-51 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W777 N$1554 N$1553 "Straight Waveguide" sch_x=-51 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W778 N$1556 N$1555 "Straight Waveguide" sch_x=-51 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W779 N$1558 N$1557 "Straight Waveguide" sch_x=-51 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W780 N$1560 N$1559 "Straight Waveguide" sch_x=-51 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W781 N$1562 N$1561 "Straight Waveguide" sch_x=-51 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W782 N$1564 N$1563 "Straight Waveguide" sch_x=-51 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W783 N$1566 N$1565 "Straight Waveguide" sch_x=-51 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W784 N$1568 N$1567 "Straight Waveguide" sch_x=-51 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W785 N$1570 N$1569 "Straight Waveguide" sch_x=-51 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W786 N$1572 N$1571 "Straight Waveguide" sch_x=-51 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W787 N$1574 N$1573 "Straight Waveguide" sch_x=-51 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W788 N$1576 N$1575 "Straight Waveguide" sch_x=-51 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W789 N$1578 N$1577 "Straight Waveguide" sch_x=-51 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W790 N$1580 N$1579 "Straight Waveguide" sch_x=-51 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W791 N$1582 N$1581 "Straight Waveguide" sch_x=-49 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W792 N$1584 N$1583 "Straight Waveguide" sch_x=-49 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W793 N$1586 N$1585 "Straight Waveguide" sch_x=-49 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W794 N$1588 N$1587 "Straight Waveguide" sch_x=-49 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W795 N$1590 N$1589 "Straight Waveguide" sch_x=-49 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W796 N$1592 N$1591 "Straight Waveguide" sch_x=-49 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W797 N$1594 N$1593 "Straight Waveguide" sch_x=-49 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W798 N$1596 N$1595 "Straight Waveguide" sch_x=-49 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W799 N$1598 N$1597 "Straight Waveguide" sch_x=-49 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W800 N$1600 N$1599 "Straight Waveguide" sch_x=-49 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W801 N$1602 N$1601 "Straight Waveguide" sch_x=-49 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W802 N$1604 N$1603 "Straight Waveguide" sch_x=-49 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W803 N$1606 N$1605 "Straight Waveguide" sch_x=-49 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W804 N$1608 N$1607 "Straight Waveguide" sch_x=-49 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W805 N$1610 N$1609 "Straight Waveguide" sch_x=-49 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W806 N$1612 N$1611 "Straight Waveguide" sch_x=-49 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W807 N$1614 N$1613 "Straight Waveguide" sch_x=-49 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W808 N$1616 N$1615 "Straight Waveguide" sch_x=-49 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W809 N$1618 N$1617 "Straight Waveguide" sch_x=-47 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W810 N$1620 N$1619 "Straight Waveguide" sch_x=-47 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W811 N$1622 N$1621 "Straight Waveguide" sch_x=-47 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W812 N$1624 N$1623 "Straight Waveguide" sch_x=-47 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W813 N$1626 N$1625 "Straight Waveguide" sch_x=-47 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W814 N$1628 N$1627 "Straight Waveguide" sch_x=-47 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W815 N$1630 N$1629 "Straight Waveguide" sch_x=-47 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W816 N$1632 N$1631 "Straight Waveguide" sch_x=-47 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W817 N$1634 N$1633 "Straight Waveguide" sch_x=-47 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W818 N$1636 N$1635 "Straight Waveguide" sch_x=-47 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W819 N$1638 N$1637 "Straight Waveguide" sch_x=-47 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W820 N$1640 N$1639 "Straight Waveguide" sch_x=-47 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W821 N$1642 N$1641 "Straight Waveguide" sch_x=-47 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W822 N$1644 N$1643 "Straight Waveguide" sch_x=-47 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W823 N$1646 N$1645 "Straight Waveguide" sch_x=-47 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W824 N$1648 N$1647 "Straight Waveguide" sch_x=-47 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W825 N$1650 N$1649 "Straight Waveguide" sch_x=-45 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W826 N$1652 N$1651 "Straight Waveguide" sch_x=-45 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W827 N$1654 N$1653 "Straight Waveguide" sch_x=-45 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W828 N$1656 N$1655 "Straight Waveguide" sch_x=-45 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W829 N$1658 N$1657 "Straight Waveguide" sch_x=-45 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W830 N$1660 N$1659 "Straight Waveguide" sch_x=-45 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W831 N$1662 N$1661 "Straight Waveguide" sch_x=-45 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W832 N$1664 N$1663 "Straight Waveguide" sch_x=-45 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W833 N$1666 N$1665 "Straight Waveguide" sch_x=-45 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W834 N$1668 N$1667 "Straight Waveguide" sch_x=-45 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W835 N$1670 N$1669 "Straight Waveguide" sch_x=-45 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W836 N$1672 N$1671 "Straight Waveguide" sch_x=-45 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W837 N$1674 N$1673 "Straight Waveguide" sch_x=-45 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W838 N$1676 N$1675 "Straight Waveguide" sch_x=-45 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W839 N$1678 N$1677 "Straight Waveguide" sch_x=-43 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W840 N$1680 N$1679 "Straight Waveguide" sch_x=-43 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W841 N$1682 N$1681 "Straight Waveguide" sch_x=-43 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W842 N$1684 N$1683 "Straight Waveguide" sch_x=-43 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W843 N$1686 N$1685 "Straight Waveguide" sch_x=-43 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W844 N$1688 N$1687 "Straight Waveguide" sch_x=-43 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W845 N$1690 N$1689 "Straight Waveguide" sch_x=-43 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W846 N$1692 N$1691 "Straight Waveguide" sch_x=-43 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W847 N$1694 N$1693 "Straight Waveguide" sch_x=-43 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W848 N$1696 N$1695 "Straight Waveguide" sch_x=-43 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W849 N$1698 N$1697 "Straight Waveguide" sch_x=-43 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W850 N$1700 N$1699 "Straight Waveguide" sch_x=-43 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W851 N$1702 N$1701 "Straight Waveguide" sch_x=-41 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W852 N$1704 N$1703 "Straight Waveguide" sch_x=-41 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W853 N$1706 N$1705 "Straight Waveguide" sch_x=-41 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W854 N$1708 N$1707 "Straight Waveguide" sch_x=-41 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W855 N$1710 N$1709 "Straight Waveguide" sch_x=-41 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W856 N$1712 N$1711 "Straight Waveguide" sch_x=-41 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W857 N$1714 N$1713 "Straight Waveguide" sch_x=-41 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W858 N$1716 N$1715 "Straight Waveguide" sch_x=-41 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W859 N$1718 N$1717 "Straight Waveguide" sch_x=-41 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W860 N$1720 N$1719 "Straight Waveguide" sch_x=-41 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W861 N$1722 N$1721 "Straight Waveguide" sch_x=-39 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W862 N$1724 N$1723 "Straight Waveguide" sch_x=-39 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W863 N$1726 N$1725 "Straight Waveguide" sch_x=-39 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W864 N$1728 N$1727 "Straight Waveguide" sch_x=-39 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W865 N$1730 N$1729 "Straight Waveguide" sch_x=-39 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W866 N$1732 N$1731 "Straight Waveguide" sch_x=-39 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W867 N$1734 N$1733 "Straight Waveguide" sch_x=-39 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W868 N$1736 N$1735 "Straight Waveguide" sch_x=-39 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W869 N$1738 N$1737 "Straight Waveguide" sch_x=-37 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W870 N$1740 N$1739 "Straight Waveguide" sch_x=-37 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W871 N$1742 N$1741 "Straight Waveguide" sch_x=-37 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W872 N$1744 N$1743 "Straight Waveguide" sch_x=-37 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W873 N$1746 N$1745 "Straight Waveguide" sch_x=-37 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W874 N$1748 N$1747 "Straight Waveguide" sch_x=-37 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W875 N$1750 N$1749 "Straight Waveguide" sch_x=-35 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W876 N$1752 N$1751 "Straight Waveguide" sch_x=-35 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W877 N$1754 N$1753 "Straight Waveguide" sch_x=-35 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W878 N$1756 N$1755 "Straight Waveguide" sch_x=-35 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W879 N$1758 N$1757 "Straight Waveguide" sch_x=-33 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W880 N$1760 N$1759 "Straight Waveguide" sch_x=-33 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W881 N$1761 N$1762 "Straight Waveguide" sch_x=-45 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W882 N$1763 N$1764 "Straight Waveguide" sch_x=-44 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W883 N$1765 N$1766 "Straight Waveguide" sch_x=-43 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W884 N$1767 N$1768 "Straight Waveguide" sch_x=-42 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W885 N$1769 N$1770 "Straight Waveguide" sch_x=-41 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W886 N$1771 N$1772 "Straight Waveguide" sch_x=-40 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W887 N$1773 N$1774 "Straight Waveguide" sch_x=-39 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W888 N$1775 N$1776 "Straight Waveguide" sch_x=-38 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W889 N$1777 N$1778 "Straight Waveguide" sch_x=-37 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W890 N$1779 N$1780 "Straight Waveguide" sch_x=-36 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W891 N$1781 N$1782 "Straight Waveguide" sch_x=-35 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W892 N$1783 N$1784 "Straight Waveguide" sch_x=-34 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W893 N$1785 N$1786 "Straight Waveguide" sch_x=-33 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W894 N$1787 N$1788 "Straight Waveguide" sch_x=-32 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W895 N$1789 N$1790 "Straight Waveguide" sch_x=-31 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W896 N$1791 N$1792 "Straight Waveguide" sch_x=-31 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W897 N$1793 N$1794 "Straight Waveguide" sch_x=-32 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W898 N$1795 N$1796 "Straight Waveguide" sch_x=-33 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W899 N$1797 N$1798 "Straight Waveguide" sch_x=-34 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W900 N$1799 N$1800 "Straight Waveguide" sch_x=-35 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W901 N$1801 N$1802 "Straight Waveguide" sch_x=-36 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W902 N$1803 N$1804 "Straight Waveguide" sch_x=-37 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W903 N$1805 N$1806 "Straight Waveguide" sch_x=-38 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W904 N$1807 N$1808 "Straight Waveguide" sch_x=-39 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W905 N$1809 N$1810 "Straight Waveguide" sch_x=-40 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W906 N$1811 N$1812 "Straight Waveguide" sch_x=-41 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W907 N$1813 N$1814 "Straight Waveguide" sch_x=-42 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W908 N$1815 N$1816 "Straight Waveguide" sch_x=-43 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W909 N$1817 N$1818 "Straight Waveguide" sch_x=-44 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W910 N$1819 N$1820 "Straight Waveguide" sch_x=-45 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W911 N$1821 N$1822 "Straight Waveguide" sch_x=-46 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W912 N$1823 N$1824 "Straight Waveguide" sch_x=-46 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W913 N$1825 N$1826 "Straight Waveguide" sch_x=61 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W914 N$1827 N$1828 "Straight Waveguide" sch_x=61 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W915 N$1829 N$1830 "Straight Waveguide" sch_x=61 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W916 N$1831 N$1832 "Straight Waveguide" sch_x=61 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W917 N$1833 N$1834 "Straight Waveguide" sch_x=61 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W918 N$1835 N$1836 "Straight Waveguide" sch_x=61 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W919 N$1837 N$1838 "Straight Waveguide" sch_x=61 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W920 N$1839 N$1840 "Straight Waveguide" sch_x=61 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W921 N$1841 N$1842 "Straight Waveguide" sch_x=61 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W922 N$1843 N$1844 "Straight Waveguide" sch_x=61 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W923 N$1845 N$1846 "Straight Waveguide" sch_x=61 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W924 N$1847 N$1848 "Straight Waveguide" sch_x=61 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W925 N$1849 N$1850 "Straight Waveguide" sch_x=61 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W926 N$1851 N$1852 "Straight Waveguide" sch_x=61 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W927 N$1853 N$1854 "Straight Waveguide" sch_x=61 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W928 N$1855 N$1856 "Straight Waveguide" sch_x=61 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W929 N$1857 N$1858 "Straight Waveguide" sch_x=61 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W930 N$1859 N$1860 "Straight Waveguide" sch_x=61 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W931 N$1861 N$1862 "Straight Waveguide" sch_x=61 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W932 N$1863 N$1864 "Straight Waveguide" sch_x=61 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W933 N$1865 N$1866 "Straight Waveguide" sch_x=61 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W934 N$1867 N$1868 "Straight Waveguide" sch_x=61 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W935 N$1869 N$1870 "Straight Waveguide" sch_x=61 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W936 N$1871 N$1872 "Straight Waveguide" sch_x=61 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W937 N$1873 N$1874 "Straight Waveguide" sch_x=61 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W938 N$1875 N$1876 "Straight Waveguide" sch_x=61 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W939 N$1877 N$1878 "Straight Waveguide" sch_x=61 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W940 N$1879 N$1880 "Straight Waveguide" sch_x=61 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W941 N$1881 N$1882 "Straight Waveguide" sch_x=61 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W942 N$1883 N$1884 "Straight Waveguide" sch_x=61 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W943 N$1885 N$1886 "Straight Waveguide" sch_x=59 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W944 N$1887 N$1888 "Straight Waveguide" sch_x=59 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W945 N$1889 N$1890 "Straight Waveguide" sch_x=59 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W946 N$1891 N$1892 "Straight Waveguide" sch_x=59 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W947 N$1893 N$1894 "Straight Waveguide" sch_x=59 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W948 N$1895 N$1896 "Straight Waveguide" sch_x=59 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W949 N$1897 N$1898 "Straight Waveguide" sch_x=59 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W950 N$1899 N$1900 "Straight Waveguide" sch_x=59 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W951 N$1901 N$1902 "Straight Waveguide" sch_x=59 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W952 N$1903 N$1904 "Straight Waveguide" sch_x=59 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W953 N$1905 N$1906 "Straight Waveguide" sch_x=59 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W954 N$1907 N$1908 "Straight Waveguide" sch_x=59 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W955 N$1909 N$1910 "Straight Waveguide" sch_x=59 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W956 N$1911 N$1912 "Straight Waveguide" sch_x=59 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W957 N$1913 N$1914 "Straight Waveguide" sch_x=59 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W958 N$1915 N$1916 "Straight Waveguide" sch_x=59 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W959 N$1917 N$1918 "Straight Waveguide" sch_x=59 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W960 N$1919 N$1920 "Straight Waveguide" sch_x=59 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W961 N$1921 N$1922 "Straight Waveguide" sch_x=59 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W962 N$1923 N$1924 "Straight Waveguide" sch_x=59 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W963 N$1925 N$1926 "Straight Waveguide" sch_x=59 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W964 N$1927 N$1928 "Straight Waveguide" sch_x=59 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W965 N$1929 N$1930 "Straight Waveguide" sch_x=59 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W966 N$1931 N$1932 "Straight Waveguide" sch_x=59 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W967 N$1933 N$1934 "Straight Waveguide" sch_x=59 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W968 N$1935 N$1936 "Straight Waveguide" sch_x=59 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W969 N$1937 N$1938 "Straight Waveguide" sch_x=59 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W970 N$1939 N$1940 "Straight Waveguide" sch_x=59 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W971 N$1941 N$1942 "Straight Waveguide" sch_x=57 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W972 N$1943 N$1944 "Straight Waveguide" sch_x=57 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W973 N$1945 N$1946 "Straight Waveguide" sch_x=57 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W974 N$1947 N$1948 "Straight Waveguide" sch_x=57 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W975 N$1949 N$1950 "Straight Waveguide" sch_x=57 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W976 N$1951 N$1952 "Straight Waveguide" sch_x=57 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W977 N$1953 N$1954 "Straight Waveguide" sch_x=57 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W978 N$1955 N$1956 "Straight Waveguide" sch_x=57 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W979 N$1957 N$1958 "Straight Waveguide" sch_x=57 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W980 N$1959 N$1960 "Straight Waveguide" sch_x=57 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W981 N$1961 N$1962 "Straight Waveguide" sch_x=57 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W982 N$1963 N$1964 "Straight Waveguide" sch_x=57 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W983 N$1965 N$1966 "Straight Waveguide" sch_x=57 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W984 N$1967 N$1968 "Straight Waveguide" sch_x=57 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W985 N$1969 N$1970 "Straight Waveguide" sch_x=57 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W986 N$1971 N$1972 "Straight Waveguide" sch_x=57 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W987 N$1973 N$1974 "Straight Waveguide" sch_x=57 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W988 N$1975 N$1976 "Straight Waveguide" sch_x=57 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W989 N$1977 N$1978 "Straight Waveguide" sch_x=57 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W990 N$1979 N$1980 "Straight Waveguide" sch_x=57 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W991 N$1981 N$1982 "Straight Waveguide" sch_x=57 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W992 N$1983 N$1984 "Straight Waveguide" sch_x=57 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W993 N$1985 N$1986 "Straight Waveguide" sch_x=57 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W994 N$1987 N$1988 "Straight Waveguide" sch_x=57 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W995 N$1989 N$1990 "Straight Waveguide" sch_x=57 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W996 N$1991 N$1992 "Straight Waveguide" sch_x=57 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W997 N$1993 N$1994 "Straight Waveguide" sch_x=55 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W998 N$1995 N$1996 "Straight Waveguide" sch_x=55 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W999 N$1997 N$1998 "Straight Waveguide" sch_x=55 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1000 N$1999 N$2000 "Straight Waveguide" sch_x=55 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1001 N$2001 N$2002 "Straight Waveguide" sch_x=55 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1002 N$2003 N$2004 "Straight Waveguide" sch_x=55 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1003 N$2005 N$2006 "Straight Waveguide" sch_x=55 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1004 N$2007 N$2008 "Straight Waveguide" sch_x=55 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1005 N$2009 N$2010 "Straight Waveguide" sch_x=55 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1006 N$2011 N$2012 "Straight Waveguide" sch_x=55 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1007 N$2013 N$2014 "Straight Waveguide" sch_x=55 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1008 N$2015 N$2016 "Straight Waveguide" sch_x=55 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1009 N$2017 N$2018 "Straight Waveguide" sch_x=55 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1010 N$2019 N$2020 "Straight Waveguide" sch_x=55 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1011 N$2021 N$2022 "Straight Waveguide" sch_x=55 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1012 N$2023 N$2024 "Straight Waveguide" sch_x=55 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1013 N$2025 N$2026 "Straight Waveguide" sch_x=55 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1014 N$2027 N$2028 "Straight Waveguide" sch_x=55 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1015 N$2029 N$2030 "Straight Waveguide" sch_x=55 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1016 N$2031 N$2032 "Straight Waveguide" sch_x=55 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1017 N$2033 N$2034 "Straight Waveguide" sch_x=55 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1018 N$2035 N$2036 "Straight Waveguide" sch_x=55 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1019 N$2037 N$2038 "Straight Waveguide" sch_x=55 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1020 N$2039 N$2040 "Straight Waveguide" sch_x=55 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1021 N$2041 N$2042 "Straight Waveguide" sch_x=53 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1022 N$2043 N$2044 "Straight Waveguide" sch_x=53 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1023 N$2045 N$2046 "Straight Waveguide" sch_x=53 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1024 N$2047 N$2048 "Straight Waveguide" sch_x=53 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1025 N$2049 N$2050 "Straight Waveguide" sch_x=53 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1026 N$2051 N$2052 "Straight Waveguide" sch_x=53 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1027 N$2053 N$2054 "Straight Waveguide" sch_x=53 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1028 N$2055 N$2056 "Straight Waveguide" sch_x=53 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1029 N$2057 N$2058 "Straight Waveguide" sch_x=53 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1030 N$2059 N$2060 "Straight Waveguide" sch_x=53 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1031 N$2061 N$2062 "Straight Waveguide" sch_x=53 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1032 N$2063 N$2064 "Straight Waveguide" sch_x=53 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1033 N$2065 N$2066 "Straight Waveguide" sch_x=53 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1034 N$2067 N$2068 "Straight Waveguide" sch_x=53 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1035 N$2069 N$2070 "Straight Waveguide" sch_x=53 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1036 N$2071 N$2072 "Straight Waveguide" sch_x=53 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1037 N$2073 N$2074 "Straight Waveguide" sch_x=53 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1038 N$2075 N$2076 "Straight Waveguide" sch_x=53 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1039 N$2077 N$2078 "Straight Waveguide" sch_x=53 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1040 N$2079 N$2080 "Straight Waveguide" sch_x=53 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1041 N$2081 N$2082 "Straight Waveguide" sch_x=53 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1042 N$2083 N$2084 "Straight Waveguide" sch_x=53 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1043 N$2085 N$2086 "Straight Waveguide" sch_x=51 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1044 N$2087 N$2088 "Straight Waveguide" sch_x=51 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1045 N$2089 N$2090 "Straight Waveguide" sch_x=51 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1046 N$2091 N$2092 "Straight Waveguide" sch_x=51 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1047 N$2093 N$2094 "Straight Waveguide" sch_x=51 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1048 N$2095 N$2096 "Straight Waveguide" sch_x=51 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1049 N$2097 N$2098 "Straight Waveguide" sch_x=51 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1050 N$2099 N$2100 "Straight Waveguide" sch_x=51 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1051 N$2101 N$2102 "Straight Waveguide" sch_x=51 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1052 N$2103 N$2104 "Straight Waveguide" sch_x=51 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1053 N$2105 N$2106 "Straight Waveguide" sch_x=51 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1054 N$2107 N$2108 "Straight Waveguide" sch_x=51 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1055 N$2109 N$2110 "Straight Waveguide" sch_x=51 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1056 N$2111 N$2112 "Straight Waveguide" sch_x=51 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1057 N$2113 N$2114 "Straight Waveguide" sch_x=51 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1058 N$2115 N$2116 "Straight Waveguide" sch_x=51 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1059 N$2117 N$2118 "Straight Waveguide" sch_x=51 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1060 N$2119 N$2120 "Straight Waveguide" sch_x=51 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1061 N$2121 N$2122 "Straight Waveguide" sch_x=51 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1062 N$2123 N$2124 "Straight Waveguide" sch_x=51 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1063 N$2125 N$2126 "Straight Waveguide" sch_x=49 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1064 N$2127 N$2128 "Straight Waveguide" sch_x=49 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1065 N$2129 N$2130 "Straight Waveguide" sch_x=49 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1066 N$2131 N$2132 "Straight Waveguide" sch_x=49 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1067 N$2133 N$2134 "Straight Waveguide" sch_x=49 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1068 N$2135 N$2136 "Straight Waveguide" sch_x=49 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1069 N$2137 N$2138 "Straight Waveguide" sch_x=49 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1070 N$2139 N$2140 "Straight Waveguide" sch_x=49 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1071 N$2141 N$2142 "Straight Waveguide" sch_x=49 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1072 N$2143 N$2144 "Straight Waveguide" sch_x=49 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1073 N$2145 N$2146 "Straight Waveguide" sch_x=49 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1074 N$2147 N$2148 "Straight Waveguide" sch_x=49 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1075 N$2149 N$2150 "Straight Waveguide" sch_x=49 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1076 N$2151 N$2152 "Straight Waveguide" sch_x=49 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1077 N$2153 N$2154 "Straight Waveguide" sch_x=49 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1078 N$2155 N$2156 "Straight Waveguide" sch_x=49 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1079 N$2157 N$2158 "Straight Waveguide" sch_x=49 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1080 N$2159 N$2160 "Straight Waveguide" sch_x=49 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1081 N$2161 N$2162 "Straight Waveguide" sch_x=47 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1082 N$2163 N$2164 "Straight Waveguide" sch_x=47 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1083 N$2165 N$2166 "Straight Waveguide" sch_x=47 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1084 N$2167 N$2168 "Straight Waveguide" sch_x=47 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1085 N$2169 N$2170 "Straight Waveguide" sch_x=47 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1086 N$2171 N$2172 "Straight Waveguide" sch_x=47 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1087 N$2173 N$2174 "Straight Waveguide" sch_x=47 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1088 N$2175 N$2176 "Straight Waveguide" sch_x=47 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1089 N$2177 N$2178 "Straight Waveguide" sch_x=47 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1090 N$2179 N$2180 "Straight Waveguide" sch_x=47 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1091 N$2181 N$2182 "Straight Waveguide" sch_x=47 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1092 N$2183 N$2184 "Straight Waveguide" sch_x=47 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1093 N$2185 N$2186 "Straight Waveguide" sch_x=47 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1094 N$2187 N$2188 "Straight Waveguide" sch_x=47 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1095 N$2189 N$2190 "Straight Waveguide" sch_x=47 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1096 N$2191 N$2192 "Straight Waveguide" sch_x=47 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1097 N$2193 N$2194 "Straight Waveguide" sch_x=45 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1098 N$2195 N$2196 "Straight Waveguide" sch_x=45 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1099 N$2197 N$2198 "Straight Waveguide" sch_x=45 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1100 N$2199 N$2200 "Straight Waveguide" sch_x=45 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1101 N$2201 N$2202 "Straight Waveguide" sch_x=45 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1102 N$2203 N$2204 "Straight Waveguide" sch_x=45 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1103 N$2205 N$2206 "Straight Waveguide" sch_x=45 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1104 N$2207 N$2208 "Straight Waveguide" sch_x=45 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1105 N$2209 N$2210 "Straight Waveguide" sch_x=45 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1106 N$2211 N$2212 "Straight Waveguide" sch_x=45 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1107 N$2213 N$2214 "Straight Waveguide" sch_x=45 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1108 N$2215 N$2216 "Straight Waveguide" sch_x=45 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1109 N$2217 N$2218 "Straight Waveguide" sch_x=45 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1110 N$2219 N$2220 "Straight Waveguide" sch_x=45 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1111 N$2221 N$2222 "Straight Waveguide" sch_x=43 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1112 N$2223 N$2224 "Straight Waveguide" sch_x=43 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1113 N$2225 N$2226 "Straight Waveguide" sch_x=43 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1114 N$2227 N$2228 "Straight Waveguide" sch_x=43 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1115 N$2229 N$2230 "Straight Waveguide" sch_x=43 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1116 N$2231 N$2232 "Straight Waveguide" sch_x=43 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1117 N$2233 N$2234 "Straight Waveguide" sch_x=43 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1118 N$2235 N$2236 "Straight Waveguide" sch_x=43 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1119 N$2237 N$2238 "Straight Waveguide" sch_x=43 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1120 N$2239 N$2240 "Straight Waveguide" sch_x=43 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1121 N$2241 N$2242 "Straight Waveguide" sch_x=43 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1122 N$2243 N$2244 "Straight Waveguide" sch_x=43 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1123 N$2245 N$2246 "Straight Waveguide" sch_x=41 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1124 N$2247 N$2248 "Straight Waveguide" sch_x=41 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1125 N$2249 N$2250 "Straight Waveguide" sch_x=41 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1126 N$2251 N$2252 "Straight Waveguide" sch_x=41 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1127 N$2253 N$2254 "Straight Waveguide" sch_x=41 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1128 N$2255 N$2256 "Straight Waveguide" sch_x=41 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1129 N$2257 N$2258 "Straight Waveguide" sch_x=41 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1130 N$2259 N$2260 "Straight Waveguide" sch_x=41 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1131 N$2261 N$2262 "Straight Waveguide" sch_x=41 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1132 N$2263 N$2264 "Straight Waveguide" sch_x=41 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1133 N$2265 N$2266 "Straight Waveguide" sch_x=39 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1134 N$2267 N$2268 "Straight Waveguide" sch_x=39 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1135 N$2269 N$2270 "Straight Waveguide" sch_x=39 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1136 N$2271 N$2272 "Straight Waveguide" sch_x=39 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1137 N$2273 N$2274 "Straight Waveguide" sch_x=39 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1138 N$2275 N$2276 "Straight Waveguide" sch_x=39 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1139 N$2277 N$2278 "Straight Waveguide" sch_x=39 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1140 N$2279 N$2280 "Straight Waveguide" sch_x=39 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1141 N$2281 N$2282 "Straight Waveguide" sch_x=37 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1142 N$2283 N$2284 "Straight Waveguide" sch_x=37 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1143 N$2285 N$2286 "Straight Waveguide" sch_x=37 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1144 N$2287 N$2288 "Straight Waveguide" sch_x=37 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1145 N$2289 N$2290 "Straight Waveguide" sch_x=37 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1146 N$2291 N$2292 "Straight Waveguide" sch_x=37 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1147 N$2293 N$2294 "Straight Waveguide" sch_x=35 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1148 N$2295 N$2296 "Straight Waveguide" sch_x=35 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1149 N$2297 N$2298 "Straight Waveguide" sch_x=35 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1150 N$2299 N$2300 "Straight Waveguide" sch_x=35 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1151 N$2301 N$2302 "Straight Waveguide" sch_x=33 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1152 N$2303 N$2304 "Straight Waveguide" sch_x=33 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1153 N$2306 N$2305 "Straight Waveguide" sch_x=45 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1154 N$2308 N$2307 "Straight Waveguide" sch_x=44 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1155 N$2310 N$2309 "Straight Waveguide" sch_x=43 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1156 N$2312 N$2311 "Straight Waveguide" sch_x=42 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1157 N$2314 N$2313 "Straight Waveguide" sch_x=41 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1158 N$2316 N$2315 "Straight Waveguide" sch_x=40 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1159 N$2318 N$2317 "Straight Waveguide" sch_x=39 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1160 N$2320 N$2319 "Straight Waveguide" sch_x=38 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1161 N$2322 N$2321 "Straight Waveguide" sch_x=37 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1162 N$2324 N$2323 "Straight Waveguide" sch_x=36 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1163 N$2326 N$2325 "Straight Waveguide" sch_x=35 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1164 N$2328 N$2327 "Straight Waveguide" sch_x=34 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1165 N$2330 N$2329 "Straight Waveguide" sch_x=33 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1166 N$2332 N$2331 "Straight Waveguide" sch_x=32 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1167 N$2334 N$2333 "Straight Waveguide" sch_x=31 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1168 N$2336 N$2335 "Straight Waveguide" sch_x=31 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1169 N$2338 N$2337 "Straight Waveguide" sch_x=32 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1170 N$2340 N$2339 "Straight Waveguide" sch_x=33 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1171 N$2342 N$2341 "Straight Waveguide" sch_x=34 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1172 N$2344 N$2343 "Straight Waveguide" sch_x=35 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1173 N$2346 N$2345 "Straight Waveguide" sch_x=36 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1174 N$2348 N$2347 "Straight Waveguide" sch_x=37 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1175 N$2350 N$2349 "Straight Waveguide" sch_x=38 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1176 N$2352 N$2351 "Straight Waveguide" sch_x=39 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1177 N$2354 N$2353 "Straight Waveguide" sch_x=40 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1178 N$2356 N$2355 "Straight Waveguide" sch_x=41 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1179 N$2358 N$2357 "Straight Waveguide" sch_x=42 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1180 N$2360 N$2359 "Straight Waveguide" sch_x=43 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1181 N$2362 N$2361 "Straight Waveguide" sch_x=44 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1182 N$2364 N$2363 "Straight Waveguide" sch_x=45 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1183 N$2366 N$2365 "Straight Waveguide" sch_x=46 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1184 N$2368 N$2367 "Straight Waveguide" sch_x=46 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1185 N$2369 N$2370 "Straight Waveguide" sch_x=-4 sch_y=-0.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1186 N$2371 N$2372 "Straight Waveguide" sch_x=-5 sch_y=-1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1187 N$2373 N$2374 "Straight Waveguide" sch_x=-5 sch_y=-2.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1188 N$2375 N$2376 "Straight Waveguide" sch_x=-3 sch_y=-1.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1189 N$2377 N$2378 "Straight Waveguide" sch_x=-3 sch_y=-2.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1190 N$2379 N$2380 "Straight Waveguide" sch_x=-4 sch_y=-3.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1191 N$2381 N$2382 "Straight Waveguide" sch_x=0 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1192 N$2383 N$2384 "Straight Waveguide" sch_x=-1 sch_y=-0.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1193 N$2385 N$2386 "Straight Waveguide" sch_x=-1 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1194 N$2387 N$2388 "Straight Waveguide" sch_x=1 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1195 N$2389 N$2390 "Straight Waveguide" sch_x=1 sch_y=-0.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1196 N$2391 N$2392 "Straight Waveguide" sch_x=0 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1197 N$2393 N$2394 "Straight Waveguide" sch_x=0 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1198 N$2395 N$2396 "Straight Waveguide" sch_x=-1 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1199 N$2397 N$2398 "Straight Waveguide" sch_x=-1 sch_y=-3.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1200 N$2399 N$2400 "Straight Waveguide" sch_x=1 sch_y=-3.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1201 N$2401 N$2402 "Straight Waveguide" sch_x=1 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1202 N$2403 N$2404 "Straight Waveguide" sch_x=0 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1203 N$2405 N$2406 "Straight Waveguide" sch_x=4 sch_y=-0.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1204 N$2407 N$2408 "Straight Waveguide" sch_x=3 sch_y=-1.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1205 N$2409 N$2410 "Straight Waveguide" sch_x=3 sch_y=-2.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1206 N$2411 N$2412 "Straight Waveguide" sch_x=5 sch_y=-2.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1207 N$2413 N$2414 "Straight Waveguide" sch_x=5 sch_y=-1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1208 N$2415 N$2416 "Straight Waveguide" sch_x=4 sch_y=-3.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1209 N$2417 N$2418 "Straight Waveguide" sch_x=-4 sch_y=-4.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1210 N$2419 N$2420 "Straight Waveguide" sch_x=-5 sch_y=-5.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1211 N$2421 N$2422 "Straight Waveguide" sch_x=-5 sch_y=-6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1212 N$2423 N$2424 "Straight Waveguide" sch_x=-3 sch_y=-5.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1213 N$2425 N$2426 "Straight Waveguide" sch_x=-3 sch_y=-6.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1214 N$2427 N$2428 "Straight Waveguide" sch_x=-4 sch_y=-7.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1215 N$2429 N$2430 "Straight Waveguide" sch_x=0 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1216 N$2431 N$2432 "Straight Waveguide" sch_x=-1 sch_y=-4.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1217 N$2433 N$2434 "Straight Waveguide" sch_x=-1 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1218 N$2435 N$2436 "Straight Waveguide" sch_x=1 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1219 N$2437 N$2438 "Straight Waveguide" sch_x=1 sch_y=-4.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1220 N$2439 N$2440 "Straight Waveguide" sch_x=0 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1221 N$2441 N$2442 "Straight Waveguide" sch_x=0 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1222 N$2443 N$2444 "Straight Waveguide" sch_x=-1 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1223 N$2445 N$2446 "Straight Waveguide" sch_x=-1 sch_y=-7.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1224 N$2447 N$2448 "Straight Waveguide" sch_x=1 sch_y=-7.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1225 N$2449 N$2450 "Straight Waveguide" sch_x=1 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1226 N$2451 N$2452 "Straight Waveguide" sch_x=0 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1227 N$2453 N$2454 "Straight Waveguide" sch_x=4 sch_y=-4.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1228 N$2455 N$2456 "Straight Waveguide" sch_x=3 sch_y=-5.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1229 N$2457 N$2458 "Straight Waveguide" sch_x=3 sch_y=-6.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1230 N$2459 N$2460 "Straight Waveguide" sch_x=5 sch_y=-6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1231 N$2461 N$2462 "Straight Waveguide" sch_x=5 sch_y=-5.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1232 N$2463 N$2464 "Straight Waveguide" sch_x=4 sch_y=-7.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1233 N$2466 N$2465 "Straight Waveguide" sch_x=-13 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1234 N$2468 N$2467 "Straight Waveguide" sch_x=-13 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1235 N$2470 N$2469 "Straight Waveguide" sch_x=-13 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1236 N$2472 N$2471 "Straight Waveguide" sch_x=-13 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1237 N$2474 N$2473 "Straight Waveguide" sch_x=-13 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1238 N$2476 N$2475 "Straight Waveguide" sch_x=-13 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1239 N$2478 N$2477 "Straight Waveguide" sch_x=-11 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1240 N$2480 N$2479 "Straight Waveguide" sch_x=-11 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1241 N$2482 N$2481 "Straight Waveguide" sch_x=-11 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1242 N$2484 N$2483 "Straight Waveguide" sch_x=-11 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1243 N$2486 N$2485 "Straight Waveguide" sch_x=-9 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1244 N$2488 N$2487 "Straight Waveguide" sch_x=-9 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1245 N$2489 N$2490 "Straight Waveguide" sch_x=-9 sch_y=-1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1246 N$2491 N$2492 "Straight Waveguide" sch_x=-8 sch_y=-2.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1247 N$2493 N$2494 "Straight Waveguide" sch_x=-7 sch_y=-3.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1248 N$2495 N$2496 "Straight Waveguide" sch_x=-7 sch_y=-4.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1249 N$2497 N$2498 "Straight Waveguide" sch_x=-8 sch_y=-5.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1250 N$2499 N$2500 "Straight Waveguide" sch_x=-9 sch_y=-6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1251 N$2501 N$2502 "Straight Waveguide" sch_x=-10 sch_y=-1.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1252 N$2503 N$2504 "Straight Waveguide" sch_x=-10 sch_y=-6.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1253 N$2505 N$2506 "Straight Waveguide" sch_x=13 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1254 N$2507 N$2508 "Straight Waveguide" sch_x=13 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1255 N$2509 N$2510 "Straight Waveguide" sch_x=13 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1256 N$2511 N$2512 "Straight Waveguide" sch_x=13 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1257 N$2513 N$2514 "Straight Waveguide" sch_x=13 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1258 N$2515 N$2516 "Straight Waveguide" sch_x=13 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1259 N$2517 N$2518 "Straight Waveguide" sch_x=11 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1260 N$2519 N$2520 "Straight Waveguide" sch_x=11 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1261 N$2521 N$2522 "Straight Waveguide" sch_x=11 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1262 N$2523 N$2524 "Straight Waveguide" sch_x=11 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1263 N$2525 N$2526 "Straight Waveguide" sch_x=9 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1264 N$2527 N$2528 "Straight Waveguide" sch_x=9 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1265 N$2530 N$2529 "Straight Waveguide" sch_x=9 sch_y=-1.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1266 N$2532 N$2531 "Straight Waveguide" sch_x=8 sch_y=-2.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1267 N$2534 N$2533 "Straight Waveguide" sch_x=7 sch_y=-3.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1268 N$2536 N$2535 "Straight Waveguide" sch_x=7 sch_y=-4.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1269 N$2538 N$2537 "Straight Waveguide" sch_x=8 sch_y=-5.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1270 N$2540 N$2539 "Straight Waveguide" sch_x=9 sch_y=-6.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1271 N$2542 N$2541 "Straight Waveguide" sch_x=10 sch_y=-1.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1272 N$2544 N$2543 "Straight Waveguide" sch_x=10 sch_y=-6.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1273 N$2545 N$2546 "Straight Waveguide" sch_x=-4 sch_y=-8.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1274 N$2547 N$2548 "Straight Waveguide" sch_x=-5 sch_y=-9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1275 N$2549 N$2550 "Straight Waveguide" sch_x=-5 sch_y=-10.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1276 N$2551 N$2552 "Straight Waveguide" sch_x=-3 sch_y=-9.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1277 N$2553 N$2554 "Straight Waveguide" sch_x=-3 sch_y=-10.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1278 N$2555 N$2556 "Straight Waveguide" sch_x=-4 sch_y=-11.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1279 N$2557 N$2558 "Straight Waveguide" sch_x=0 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1280 N$2559 N$2560 "Straight Waveguide" sch_x=-1 sch_y=-8.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1281 N$2561 N$2562 "Straight Waveguide" sch_x=-1 sch_y=-9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1282 N$2563 N$2564 "Straight Waveguide" sch_x=1 sch_y=-9.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1283 N$2565 N$2566 "Straight Waveguide" sch_x=1 sch_y=-8.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1284 N$2567 N$2568 "Straight Waveguide" sch_x=0 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1285 N$2569 N$2570 "Straight Waveguide" sch_x=0 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1286 N$2571 N$2572 "Straight Waveguide" sch_x=-1 sch_y=-10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1287 N$2573 N$2574 "Straight Waveguide" sch_x=-1 sch_y=-11.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1288 N$2575 N$2576 "Straight Waveguide" sch_x=1 sch_y=-11.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1289 N$2577 N$2578 "Straight Waveguide" sch_x=1 sch_y=-10.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1290 N$2579 N$2580 "Straight Waveguide" sch_x=0 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1291 N$2581 N$2582 "Straight Waveguide" sch_x=4 sch_y=-8.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1292 N$2583 N$2584 "Straight Waveguide" sch_x=3 sch_y=-9.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1293 N$2585 N$2586 "Straight Waveguide" sch_x=3 sch_y=-10.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1294 N$2587 N$2588 "Straight Waveguide" sch_x=5 sch_y=-10.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1295 N$2589 N$2590 "Straight Waveguide" sch_x=5 sch_y=-9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1296 N$2591 N$2592 "Straight Waveguide" sch_x=4 sch_y=-11.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1297 N$2593 N$2594 "Straight Waveguide" sch_x=-4 sch_y=-12.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1298 N$2595 N$2596 "Straight Waveguide" sch_x=-5 sch_y=-13.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1299 N$2597 N$2598 "Straight Waveguide" sch_x=-5 sch_y=-14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1300 N$2599 N$2600 "Straight Waveguide" sch_x=-3 sch_y=-13.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1301 N$2601 N$2602 "Straight Waveguide" sch_x=-3 sch_y=-14.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1302 N$2603 N$2604 "Straight Waveguide" sch_x=-4 sch_y=-15.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1303 N$2605 N$2606 "Straight Waveguide" sch_x=0 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1304 N$2607 N$2608 "Straight Waveguide" sch_x=-1 sch_y=-12.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1305 N$2609 N$2610 "Straight Waveguide" sch_x=-1 sch_y=-13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1306 N$2611 N$2612 "Straight Waveguide" sch_x=1 sch_y=-13.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1307 N$2613 N$2614 "Straight Waveguide" sch_x=1 sch_y=-12.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1308 N$2615 N$2616 "Straight Waveguide" sch_x=0 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1309 N$2617 N$2618 "Straight Waveguide" sch_x=0 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1310 N$2619 N$2620 "Straight Waveguide" sch_x=-1 sch_y=-14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1311 N$2621 N$2622 "Straight Waveguide" sch_x=-1 sch_y=-15.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1312 N$2623 N$2624 "Straight Waveguide" sch_x=1 sch_y=-15.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1313 N$2625 N$2626 "Straight Waveguide" sch_x=1 sch_y=-14.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1314 N$2627 N$2628 "Straight Waveguide" sch_x=0 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1315 N$2629 N$2630 "Straight Waveguide" sch_x=4 sch_y=-12.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1316 N$2631 N$2632 "Straight Waveguide" sch_x=3 sch_y=-13.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1317 N$2633 N$2634 "Straight Waveguide" sch_x=3 sch_y=-14.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1318 N$2635 N$2636 "Straight Waveguide" sch_x=5 sch_y=-14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1319 N$2637 N$2638 "Straight Waveguide" sch_x=5 sch_y=-13.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1320 N$2639 N$2640 "Straight Waveguide" sch_x=4 sch_y=-15.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1321 N$2642 N$2641 "Straight Waveguide" sch_x=-13 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1322 N$2644 N$2643 "Straight Waveguide" sch_x=-13 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1323 N$2646 N$2645 "Straight Waveguide" sch_x=-13 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1324 N$2648 N$2647 "Straight Waveguide" sch_x=-13 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1325 N$2650 N$2649 "Straight Waveguide" sch_x=-13 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1326 N$2652 N$2651 "Straight Waveguide" sch_x=-13 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1327 N$2654 N$2653 "Straight Waveguide" sch_x=-11 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1328 N$2656 N$2655 "Straight Waveguide" sch_x=-11 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1329 N$2658 N$2657 "Straight Waveguide" sch_x=-11 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1330 N$2660 N$2659 "Straight Waveguide" sch_x=-11 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1331 N$2662 N$2661 "Straight Waveguide" sch_x=-9 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1332 N$2664 N$2663 "Straight Waveguide" sch_x=-9 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1333 N$2665 N$2666 "Straight Waveguide" sch_x=-9 sch_y=-9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1334 N$2667 N$2668 "Straight Waveguide" sch_x=-8 sch_y=-10.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1335 N$2669 N$2670 "Straight Waveguide" sch_x=-7 sch_y=-11.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1336 N$2671 N$2672 "Straight Waveguide" sch_x=-7 sch_y=-12.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1337 N$2673 N$2674 "Straight Waveguide" sch_x=-8 sch_y=-13.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1338 N$2675 N$2676 "Straight Waveguide" sch_x=-9 sch_y=-14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1339 N$2677 N$2678 "Straight Waveguide" sch_x=-10 sch_y=-9.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1340 N$2679 N$2680 "Straight Waveguide" sch_x=-10 sch_y=-14.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1341 N$2681 N$2682 "Straight Waveguide" sch_x=13 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1342 N$2683 N$2684 "Straight Waveguide" sch_x=13 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1343 N$2685 N$2686 "Straight Waveguide" sch_x=13 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1344 N$2687 N$2688 "Straight Waveguide" sch_x=13 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1345 N$2689 N$2690 "Straight Waveguide" sch_x=13 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1346 N$2691 N$2692 "Straight Waveguide" sch_x=13 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1347 N$2693 N$2694 "Straight Waveguide" sch_x=11 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1348 N$2695 N$2696 "Straight Waveguide" sch_x=11 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1349 N$2697 N$2698 "Straight Waveguide" sch_x=11 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1350 N$2699 N$2700 "Straight Waveguide" sch_x=11 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1351 N$2701 N$2702 "Straight Waveguide" sch_x=9 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1352 N$2703 N$2704 "Straight Waveguide" sch_x=9 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1353 N$2706 N$2705 "Straight Waveguide" sch_x=9 sch_y=-9.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1354 N$2708 N$2707 "Straight Waveguide" sch_x=8 sch_y=-10.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1355 N$2710 N$2709 "Straight Waveguide" sch_x=7 sch_y=-11.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1356 N$2712 N$2711 "Straight Waveguide" sch_x=7 sch_y=-12.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1357 N$2714 N$2713 "Straight Waveguide" sch_x=8 sch_y=-13.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1358 N$2716 N$2715 "Straight Waveguide" sch_x=9 sch_y=-14.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1359 N$2718 N$2717 "Straight Waveguide" sch_x=10 sch_y=-9.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1360 N$2720 N$2719 "Straight Waveguide" sch_x=10 sch_y=-14.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1361 N$2722 N$2721 "Straight Waveguide" sch_x=-29 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1362 N$2724 N$2723 "Straight Waveguide" sch_x=-29 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1363 N$2726 N$2725 "Straight Waveguide" sch_x=-29 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1364 N$2728 N$2727 "Straight Waveguide" sch_x=-29 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1365 N$2730 N$2729 "Straight Waveguide" sch_x=-29 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1366 N$2732 N$2731 "Straight Waveguide" sch_x=-29 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1367 N$2734 N$2733 "Straight Waveguide" sch_x=-29 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1368 N$2736 N$2735 "Straight Waveguide" sch_x=-29 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1369 N$2738 N$2737 "Straight Waveguide" sch_x=-29 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1370 N$2740 N$2739 "Straight Waveguide" sch_x=-29 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1371 N$2742 N$2741 "Straight Waveguide" sch_x=-29 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1372 N$2744 N$2743 "Straight Waveguide" sch_x=-29 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1373 N$2746 N$2745 "Straight Waveguide" sch_x=-29 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1374 N$2748 N$2747 "Straight Waveguide" sch_x=-29 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1375 N$2750 N$2749 "Straight Waveguide" sch_x=-27 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1376 N$2752 N$2751 "Straight Waveguide" sch_x=-27 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1377 N$2754 N$2753 "Straight Waveguide" sch_x=-27 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1378 N$2756 N$2755 "Straight Waveguide" sch_x=-27 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1379 N$2758 N$2757 "Straight Waveguide" sch_x=-27 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1380 N$2760 N$2759 "Straight Waveguide" sch_x=-27 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1381 N$2762 N$2761 "Straight Waveguide" sch_x=-27 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1382 N$2764 N$2763 "Straight Waveguide" sch_x=-27 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1383 N$2766 N$2765 "Straight Waveguide" sch_x=-27 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1384 N$2768 N$2767 "Straight Waveguide" sch_x=-27 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1385 N$2770 N$2769 "Straight Waveguide" sch_x=-27 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1386 N$2772 N$2771 "Straight Waveguide" sch_x=-27 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1387 N$2774 N$2773 "Straight Waveguide" sch_x=-25 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1388 N$2776 N$2775 "Straight Waveguide" sch_x=-25 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1389 N$2778 N$2777 "Straight Waveguide" sch_x=-25 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1390 N$2780 N$2779 "Straight Waveguide" sch_x=-25 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1391 N$2782 N$2781 "Straight Waveguide" sch_x=-25 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1392 N$2784 N$2783 "Straight Waveguide" sch_x=-25 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1393 N$2786 N$2785 "Straight Waveguide" sch_x=-25 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1394 N$2788 N$2787 "Straight Waveguide" sch_x=-25 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1395 N$2790 N$2789 "Straight Waveguide" sch_x=-25 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1396 N$2792 N$2791 "Straight Waveguide" sch_x=-25 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1397 N$2794 N$2793 "Straight Waveguide" sch_x=-23 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1398 N$2796 N$2795 "Straight Waveguide" sch_x=-23 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1399 N$2798 N$2797 "Straight Waveguide" sch_x=-23 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1400 N$2800 N$2799 "Straight Waveguide" sch_x=-23 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1401 N$2802 N$2801 "Straight Waveguide" sch_x=-23 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1402 N$2804 N$2803 "Straight Waveguide" sch_x=-23 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1403 N$2806 N$2805 "Straight Waveguide" sch_x=-23 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1404 N$2808 N$2807 "Straight Waveguide" sch_x=-23 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1405 N$2810 N$2809 "Straight Waveguide" sch_x=-21 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1406 N$2812 N$2811 "Straight Waveguide" sch_x=-21 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1407 N$2814 N$2813 "Straight Waveguide" sch_x=-21 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1408 N$2816 N$2815 "Straight Waveguide" sch_x=-21 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1409 N$2818 N$2817 "Straight Waveguide" sch_x=-21 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1410 N$2820 N$2819 "Straight Waveguide" sch_x=-21 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1411 N$2822 N$2821 "Straight Waveguide" sch_x=-19 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1412 N$2824 N$2823 "Straight Waveguide" sch_x=-19 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1413 N$2826 N$2825 "Straight Waveguide" sch_x=-19 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1414 N$2828 N$2827 "Straight Waveguide" sch_x=-19 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1415 N$2830 N$2829 "Straight Waveguide" sch_x=-17 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1416 N$2832 N$2831 "Straight Waveguide" sch_x=-17 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1417 N$2833 N$2834 "Straight Waveguide" sch_x=-21 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1418 N$2835 N$2836 "Straight Waveguide" sch_x=-20 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1419 N$2837 N$2838 "Straight Waveguide" sch_x=-19 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1420 N$2839 N$2840 "Straight Waveguide" sch_x=-18 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1421 N$2841 N$2842 "Straight Waveguide" sch_x=-17 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1422 N$2843 N$2844 "Straight Waveguide" sch_x=-16 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1423 N$2845 N$2846 "Straight Waveguide" sch_x=-15 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1424 N$2847 N$2848 "Straight Waveguide" sch_x=-15 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1425 N$2849 N$2850 "Straight Waveguide" sch_x=-16 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1426 N$2851 N$2852 "Straight Waveguide" sch_x=-17 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1427 N$2853 N$2854 "Straight Waveguide" sch_x=-18 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1428 N$2855 N$2856 "Straight Waveguide" sch_x=-19 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1429 N$2857 N$2858 "Straight Waveguide" sch_x=-20 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1430 N$2859 N$2860 "Straight Waveguide" sch_x=-21 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1431 N$2861 N$2862 "Straight Waveguide" sch_x=-22 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1432 N$2863 N$2864 "Straight Waveguide" sch_x=-22 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1433 N$2865 N$2866 "Straight Waveguide" sch_x=29 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1434 N$2867 N$2868 "Straight Waveguide" sch_x=29 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1435 N$2869 N$2870 "Straight Waveguide" sch_x=29 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1436 N$2871 N$2872 "Straight Waveguide" sch_x=29 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1437 N$2873 N$2874 "Straight Waveguide" sch_x=29 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1438 N$2875 N$2876 "Straight Waveguide" sch_x=29 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1439 N$2877 N$2878 "Straight Waveguide" sch_x=29 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1440 N$2879 N$2880 "Straight Waveguide" sch_x=29 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1441 N$2881 N$2882 "Straight Waveguide" sch_x=29 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1442 N$2883 N$2884 "Straight Waveguide" sch_x=29 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1443 N$2885 N$2886 "Straight Waveguide" sch_x=29 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1444 N$2887 N$2888 "Straight Waveguide" sch_x=29 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1445 N$2889 N$2890 "Straight Waveguide" sch_x=29 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1446 N$2891 N$2892 "Straight Waveguide" sch_x=29 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1447 N$2893 N$2894 "Straight Waveguide" sch_x=27 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1448 N$2895 N$2896 "Straight Waveguide" sch_x=27 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1449 N$2897 N$2898 "Straight Waveguide" sch_x=27 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1450 N$2899 N$2900 "Straight Waveguide" sch_x=27 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1451 N$2901 N$2902 "Straight Waveguide" sch_x=27 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1452 N$2903 N$2904 "Straight Waveguide" sch_x=27 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1453 N$2905 N$2906 "Straight Waveguide" sch_x=27 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1454 N$2907 N$2908 "Straight Waveguide" sch_x=27 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1455 N$2909 N$2910 "Straight Waveguide" sch_x=27 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1456 N$2911 N$2912 "Straight Waveguide" sch_x=27 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1457 N$2913 N$2914 "Straight Waveguide" sch_x=27 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1458 N$2915 N$2916 "Straight Waveguide" sch_x=27 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1459 N$2917 N$2918 "Straight Waveguide" sch_x=25 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1460 N$2919 N$2920 "Straight Waveguide" sch_x=25 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1461 N$2921 N$2922 "Straight Waveguide" sch_x=25 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1462 N$2923 N$2924 "Straight Waveguide" sch_x=25 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1463 N$2925 N$2926 "Straight Waveguide" sch_x=25 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1464 N$2927 N$2928 "Straight Waveguide" sch_x=25 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1465 N$2929 N$2930 "Straight Waveguide" sch_x=25 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1466 N$2931 N$2932 "Straight Waveguide" sch_x=25 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1467 N$2933 N$2934 "Straight Waveguide" sch_x=25 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1468 N$2935 N$2936 "Straight Waveguide" sch_x=25 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1469 N$2937 N$2938 "Straight Waveguide" sch_x=23 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1470 N$2939 N$2940 "Straight Waveguide" sch_x=23 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1471 N$2941 N$2942 "Straight Waveguide" sch_x=23 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1472 N$2943 N$2944 "Straight Waveguide" sch_x=23 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1473 N$2945 N$2946 "Straight Waveguide" sch_x=23 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1474 N$2947 N$2948 "Straight Waveguide" sch_x=23 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1475 N$2949 N$2950 "Straight Waveguide" sch_x=23 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1476 N$2951 N$2952 "Straight Waveguide" sch_x=23 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1477 N$2953 N$2954 "Straight Waveguide" sch_x=21 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1478 N$2955 N$2956 "Straight Waveguide" sch_x=21 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1479 N$2957 N$2958 "Straight Waveguide" sch_x=21 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1480 N$2959 N$2960 "Straight Waveguide" sch_x=21 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1481 N$2961 N$2962 "Straight Waveguide" sch_x=21 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1482 N$2963 N$2964 "Straight Waveguide" sch_x=21 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1483 N$2965 N$2966 "Straight Waveguide" sch_x=19 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1484 N$2967 N$2968 "Straight Waveguide" sch_x=19 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1485 N$2969 N$2970 "Straight Waveguide" sch_x=19 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1486 N$2971 N$2972 "Straight Waveguide" sch_x=19 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1487 N$2973 N$2974 "Straight Waveguide" sch_x=17 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1488 N$2975 N$2976 "Straight Waveguide" sch_x=17 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1489 N$2978 N$2977 "Straight Waveguide" sch_x=21 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1490 N$2980 N$2979 "Straight Waveguide" sch_x=20 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1491 N$2982 N$2981 "Straight Waveguide" sch_x=19 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1492 N$2984 N$2983 "Straight Waveguide" sch_x=18 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1493 N$2986 N$2985 "Straight Waveguide" sch_x=17 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1494 N$2988 N$2987 "Straight Waveguide" sch_x=16 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1495 N$2990 N$2989 "Straight Waveguide" sch_x=15 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1496 N$2992 N$2991 "Straight Waveguide" sch_x=15 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1497 N$2994 N$2993 "Straight Waveguide" sch_x=16 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1498 N$2996 N$2995 "Straight Waveguide" sch_x=17 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1499 N$2998 N$2997 "Straight Waveguide" sch_x=18 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1500 N$3000 N$2999 "Straight Waveguide" sch_x=19 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1501 N$3002 N$3001 "Straight Waveguide" sch_x=20 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1502 N$3004 N$3003 "Straight Waveguide" sch_x=21 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1503 N$3006 N$3005 "Straight Waveguide" sch_x=22 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1504 N$3008 N$3007 "Straight Waveguide" sch_x=22 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1505 N$3009 N$3010 "Straight Waveguide" sch_x=-4 sch_y=-16.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1506 N$3011 N$3012 "Straight Waveguide" sch_x=-5 sch_y=-17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1507 N$3013 N$3014 "Straight Waveguide" sch_x=-5 sch_y=-18.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1508 N$3015 N$3016 "Straight Waveguide" sch_x=-3 sch_y=-17.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1509 N$3017 N$3018 "Straight Waveguide" sch_x=-3 sch_y=-18.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1510 N$3019 N$3020 "Straight Waveguide" sch_x=-4 sch_y=-19.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1511 N$3021 N$3022 "Straight Waveguide" sch_x=0 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1512 N$3023 N$3024 "Straight Waveguide" sch_x=-1 sch_y=-16.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1513 N$3025 N$3026 "Straight Waveguide" sch_x=-1 sch_y=-17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1514 N$3027 N$3028 "Straight Waveguide" sch_x=1 sch_y=-17.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1515 N$3029 N$3030 "Straight Waveguide" sch_x=1 sch_y=-16.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1516 N$3031 N$3032 "Straight Waveguide" sch_x=0 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1517 N$3033 N$3034 "Straight Waveguide" sch_x=0 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1518 N$3035 N$3036 "Straight Waveguide" sch_x=-1 sch_y=-18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1519 N$3037 N$3038 "Straight Waveguide" sch_x=-1 sch_y=-19.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1520 N$3039 N$3040 "Straight Waveguide" sch_x=1 sch_y=-19.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1521 N$3041 N$3042 "Straight Waveguide" sch_x=1 sch_y=-18.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1522 N$3043 N$3044 "Straight Waveguide" sch_x=0 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1523 N$3045 N$3046 "Straight Waveguide" sch_x=4 sch_y=-16.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1524 N$3047 N$3048 "Straight Waveguide" sch_x=3 sch_y=-17.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1525 N$3049 N$3050 "Straight Waveguide" sch_x=3 sch_y=-18.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1526 N$3051 N$3052 "Straight Waveguide" sch_x=5 sch_y=-18.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1527 N$3053 N$3054 "Straight Waveguide" sch_x=5 sch_y=-17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1528 N$3055 N$3056 "Straight Waveguide" sch_x=4 sch_y=-19.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1529 N$3057 N$3058 "Straight Waveguide" sch_x=-4 sch_y=-20.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1530 N$3059 N$3060 "Straight Waveguide" sch_x=-5 sch_y=-21.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1531 N$3061 N$3062 "Straight Waveguide" sch_x=-5 sch_y=-22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1532 N$3063 N$3064 "Straight Waveguide" sch_x=-3 sch_y=-21.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1533 N$3065 N$3066 "Straight Waveguide" sch_x=-3 sch_y=-22.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1534 N$3067 N$3068 "Straight Waveguide" sch_x=-4 sch_y=-23.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1535 N$3069 N$3070 "Straight Waveguide" sch_x=0 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1536 N$3071 N$3072 "Straight Waveguide" sch_x=-1 sch_y=-20.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1537 N$3073 N$3074 "Straight Waveguide" sch_x=-1 sch_y=-21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1538 N$3075 N$3076 "Straight Waveguide" sch_x=1 sch_y=-21.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1539 N$3077 N$3078 "Straight Waveguide" sch_x=1 sch_y=-20.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1540 N$3079 N$3080 "Straight Waveguide" sch_x=0 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1541 N$3081 N$3082 "Straight Waveguide" sch_x=0 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1542 N$3083 N$3084 "Straight Waveguide" sch_x=-1 sch_y=-22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1543 N$3085 N$3086 "Straight Waveguide" sch_x=-1 sch_y=-23.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1544 N$3087 N$3088 "Straight Waveguide" sch_x=1 sch_y=-23.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1545 N$3089 N$3090 "Straight Waveguide" sch_x=1 sch_y=-22.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1546 N$3091 N$3092 "Straight Waveguide" sch_x=0 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1547 N$3093 N$3094 "Straight Waveguide" sch_x=4 sch_y=-20.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1548 N$3095 N$3096 "Straight Waveguide" sch_x=3 sch_y=-21.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1549 N$3097 N$3098 "Straight Waveguide" sch_x=3 sch_y=-22.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1550 N$3099 N$3100 "Straight Waveguide" sch_x=5 sch_y=-22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1551 N$3101 N$3102 "Straight Waveguide" sch_x=5 sch_y=-21.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1552 N$3103 N$3104 "Straight Waveguide" sch_x=4 sch_y=-23.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1553 N$3106 N$3105 "Straight Waveguide" sch_x=-13 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1554 N$3108 N$3107 "Straight Waveguide" sch_x=-13 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1555 N$3110 N$3109 "Straight Waveguide" sch_x=-13 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1556 N$3112 N$3111 "Straight Waveguide" sch_x=-13 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1557 N$3114 N$3113 "Straight Waveguide" sch_x=-13 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1558 N$3116 N$3115 "Straight Waveguide" sch_x=-13 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1559 N$3118 N$3117 "Straight Waveguide" sch_x=-11 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1560 N$3120 N$3119 "Straight Waveguide" sch_x=-11 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1561 N$3122 N$3121 "Straight Waveguide" sch_x=-11 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1562 N$3124 N$3123 "Straight Waveguide" sch_x=-11 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1563 N$3126 N$3125 "Straight Waveguide" sch_x=-9 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1564 N$3128 N$3127 "Straight Waveguide" sch_x=-9 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1565 N$3129 N$3130 "Straight Waveguide" sch_x=-9 sch_y=-17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1566 N$3131 N$3132 "Straight Waveguide" sch_x=-8 sch_y=-18.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1567 N$3133 N$3134 "Straight Waveguide" sch_x=-7 sch_y=-19.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1568 N$3135 N$3136 "Straight Waveguide" sch_x=-7 sch_y=-20.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1569 N$3137 N$3138 "Straight Waveguide" sch_x=-8 sch_y=-21.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1570 N$3139 N$3140 "Straight Waveguide" sch_x=-9 sch_y=-22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1571 N$3141 N$3142 "Straight Waveguide" sch_x=-10 sch_y=-17.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1572 N$3143 N$3144 "Straight Waveguide" sch_x=-10 sch_y=-22.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1573 N$3145 N$3146 "Straight Waveguide" sch_x=13 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1574 N$3147 N$3148 "Straight Waveguide" sch_x=13 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1575 N$3149 N$3150 "Straight Waveguide" sch_x=13 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1576 N$3151 N$3152 "Straight Waveguide" sch_x=13 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1577 N$3153 N$3154 "Straight Waveguide" sch_x=13 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1578 N$3155 N$3156 "Straight Waveguide" sch_x=13 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1579 N$3157 N$3158 "Straight Waveguide" sch_x=11 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1580 N$3159 N$3160 "Straight Waveguide" sch_x=11 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1581 N$3161 N$3162 "Straight Waveguide" sch_x=11 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1582 N$3163 N$3164 "Straight Waveguide" sch_x=11 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1583 N$3165 N$3166 "Straight Waveguide" sch_x=9 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1584 N$3167 N$3168 "Straight Waveguide" sch_x=9 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1585 N$3170 N$3169 "Straight Waveguide" sch_x=9 sch_y=-17.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1586 N$3172 N$3171 "Straight Waveguide" sch_x=8 sch_y=-18.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1587 N$3174 N$3173 "Straight Waveguide" sch_x=7 sch_y=-19.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1588 N$3176 N$3175 "Straight Waveguide" sch_x=7 sch_y=-20.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1589 N$3178 N$3177 "Straight Waveguide" sch_x=8 sch_y=-21.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1590 N$3180 N$3179 "Straight Waveguide" sch_x=9 sch_y=-22.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1591 N$3182 N$3181 "Straight Waveguide" sch_x=10 sch_y=-17.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1592 N$3184 N$3183 "Straight Waveguide" sch_x=10 sch_y=-22.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1593 N$3185 N$3186 "Straight Waveguide" sch_x=-4 sch_y=-24.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1594 N$3187 N$3188 "Straight Waveguide" sch_x=-5 sch_y=-25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1595 N$3189 N$3190 "Straight Waveguide" sch_x=-5 sch_y=-26.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1596 N$3191 N$3192 "Straight Waveguide" sch_x=-3 sch_y=-25.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1597 N$3193 N$3194 "Straight Waveguide" sch_x=-3 sch_y=-26.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1598 N$3195 N$3196 "Straight Waveguide" sch_x=-4 sch_y=-27.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1599 N$3197 N$3198 "Straight Waveguide" sch_x=0 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1600 N$3199 N$3200 "Straight Waveguide" sch_x=-1 sch_y=-24.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1601 N$3201 N$3202 "Straight Waveguide" sch_x=-1 sch_y=-25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1602 N$3203 N$3204 "Straight Waveguide" sch_x=1 sch_y=-25.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1603 N$3205 N$3206 "Straight Waveguide" sch_x=1 sch_y=-24.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1604 N$3207 N$3208 "Straight Waveguide" sch_x=0 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1605 N$3209 N$3210 "Straight Waveguide" sch_x=0 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1606 N$3211 N$3212 "Straight Waveguide" sch_x=-1 sch_y=-26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1607 N$3213 N$3214 "Straight Waveguide" sch_x=-1 sch_y=-27.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1608 N$3215 N$3216 "Straight Waveguide" sch_x=1 sch_y=-27.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1609 N$3217 N$3218 "Straight Waveguide" sch_x=1 sch_y=-26.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1610 N$3219 N$3220 "Straight Waveguide" sch_x=0 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1611 N$3221 N$3222 "Straight Waveguide" sch_x=4 sch_y=-24.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1612 N$3223 N$3224 "Straight Waveguide" sch_x=3 sch_y=-25.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1613 N$3225 N$3226 "Straight Waveguide" sch_x=3 sch_y=-26.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1614 N$3227 N$3228 "Straight Waveguide" sch_x=5 sch_y=-26.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1615 N$3229 N$3230 "Straight Waveguide" sch_x=5 sch_y=-25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1616 N$3231 N$3232 "Straight Waveguide" sch_x=4 sch_y=-27.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1617 N$3233 N$3234 "Straight Waveguide" sch_x=-4 sch_y=-28.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1618 N$3235 N$3236 "Straight Waveguide" sch_x=-5 sch_y=-29.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1619 N$3237 N$3238 "Straight Waveguide" sch_x=-5 sch_y=-30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1620 N$3239 N$3240 "Straight Waveguide" sch_x=-3 sch_y=-29.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1621 N$3241 N$3242 "Straight Waveguide" sch_x=-3 sch_y=-30.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1622 N$3243 N$3244 "Straight Waveguide" sch_x=-4 sch_y=-31.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1623 N$3245 N$3246 "Straight Waveguide" sch_x=0 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1624 N$3247 N$3248 "Straight Waveguide" sch_x=-1 sch_y=-28.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1625 N$3249 N$3250 "Straight Waveguide" sch_x=-1 sch_y=-29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1626 N$3251 N$3252 "Straight Waveguide" sch_x=1 sch_y=-29.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1627 N$3253 N$3254 "Straight Waveguide" sch_x=1 sch_y=-28.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1628 N$3255 N$3256 "Straight Waveguide" sch_x=0 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1629 N$3257 N$3258 "Straight Waveguide" sch_x=0 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1630 N$3259 N$3260 "Straight Waveguide" sch_x=-1 sch_y=-30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1631 N$3261 N$3262 "Straight Waveguide" sch_x=-1 sch_y=-31.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1632 N$3263 N$3264 "Straight Waveguide" sch_x=1 sch_y=-31.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1633 N$3265 N$3266 "Straight Waveguide" sch_x=1 sch_y=-30.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1634 N$3267 N$3268 "Straight Waveguide" sch_x=0 sch_y=-31.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1635 N$3269 N$3270 "Straight Waveguide" sch_x=4 sch_y=-28.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1636 N$3271 N$3272 "Straight Waveguide" sch_x=3 sch_y=-29.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1637 N$3273 N$3274 "Straight Waveguide" sch_x=3 sch_y=-30.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1638 N$3275 N$3276 "Straight Waveguide" sch_x=5 sch_y=-30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1639 N$3277 N$3278 "Straight Waveguide" sch_x=5 sch_y=-29.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1640 N$3279 N$3280 "Straight Waveguide" sch_x=4 sch_y=-31.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1641 N$3282 N$3281 "Straight Waveguide" sch_x=-13 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1642 N$3284 N$3283 "Straight Waveguide" sch_x=-13 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1643 N$3286 N$3285 "Straight Waveguide" sch_x=-13 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1644 N$3288 N$3287 "Straight Waveguide" sch_x=-13 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1645 N$3290 N$3289 "Straight Waveguide" sch_x=-13 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1646 N$3292 N$3291 "Straight Waveguide" sch_x=-13 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1647 N$3294 N$3293 "Straight Waveguide" sch_x=-11 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1648 N$3296 N$3295 "Straight Waveguide" sch_x=-11 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1649 N$3298 N$3297 "Straight Waveguide" sch_x=-11 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1650 N$3300 N$3299 "Straight Waveguide" sch_x=-11 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1651 N$3302 N$3301 "Straight Waveguide" sch_x=-9 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1652 N$3304 N$3303 "Straight Waveguide" sch_x=-9 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1653 N$3305 N$3306 "Straight Waveguide" sch_x=-9 sch_y=-25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1654 N$3307 N$3308 "Straight Waveguide" sch_x=-8 sch_y=-26.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1655 N$3309 N$3310 "Straight Waveguide" sch_x=-7 sch_y=-27.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1656 N$3311 N$3312 "Straight Waveguide" sch_x=-7 sch_y=-28.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1657 N$3313 N$3314 "Straight Waveguide" sch_x=-8 sch_y=-29.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1658 N$3315 N$3316 "Straight Waveguide" sch_x=-9 sch_y=-30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1659 N$3317 N$3318 "Straight Waveguide" sch_x=-10 sch_y=-25.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1660 N$3319 N$3320 "Straight Waveguide" sch_x=-10 sch_y=-30.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1661 N$3321 N$3322 "Straight Waveguide" sch_x=13 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1662 N$3323 N$3324 "Straight Waveguide" sch_x=13 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1663 N$3325 N$3326 "Straight Waveguide" sch_x=13 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1664 N$3327 N$3328 "Straight Waveguide" sch_x=13 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1665 N$3329 N$3330 "Straight Waveguide" sch_x=13 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1666 N$3331 N$3332 "Straight Waveguide" sch_x=13 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1667 N$3333 N$3334 "Straight Waveguide" sch_x=11 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1668 N$3335 N$3336 "Straight Waveguide" sch_x=11 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1669 N$3337 N$3338 "Straight Waveguide" sch_x=11 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1670 N$3339 N$3340 "Straight Waveguide" sch_x=11 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1671 N$3341 N$3342 "Straight Waveguide" sch_x=9 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1672 N$3343 N$3344 "Straight Waveguide" sch_x=9 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1673 N$3346 N$3345 "Straight Waveguide" sch_x=9 sch_y=-25.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1674 N$3348 N$3347 "Straight Waveguide" sch_x=8 sch_y=-26.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1675 N$3350 N$3349 "Straight Waveguide" sch_x=7 sch_y=-27.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1676 N$3352 N$3351 "Straight Waveguide" sch_x=7 sch_y=-28.625 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1677 N$3354 N$3353 "Straight Waveguide" sch_x=8 sch_y=-29.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1678 N$3356 N$3355 "Straight Waveguide" sch_x=9 sch_y=-30.375 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1679 N$3358 N$3357 "Straight Waveguide" sch_x=10 sch_y=-25.125 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1680 N$3360 N$3359 "Straight Waveguide" sch_x=10 sch_y=-30.875 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1681 N$3362 N$3361 "Straight Waveguide" sch_x=-29 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1682 N$3364 N$3363 "Straight Waveguide" sch_x=-29 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1683 N$3366 N$3365 "Straight Waveguide" sch_x=-29 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1684 N$3368 N$3367 "Straight Waveguide" sch_x=-29 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1685 N$3370 N$3369 "Straight Waveguide" sch_x=-29 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1686 N$3372 N$3371 "Straight Waveguide" sch_x=-29 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1687 N$3374 N$3373 "Straight Waveguide" sch_x=-29 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1688 N$3376 N$3375 "Straight Waveguide" sch_x=-29 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1689 N$3378 N$3377 "Straight Waveguide" sch_x=-29 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1690 N$3380 N$3379 "Straight Waveguide" sch_x=-29 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1691 N$3382 N$3381 "Straight Waveguide" sch_x=-29 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1692 N$3384 N$3383 "Straight Waveguide" sch_x=-29 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1693 N$3386 N$3385 "Straight Waveguide" sch_x=-29 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1694 N$3388 N$3387 "Straight Waveguide" sch_x=-29 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1695 N$3390 N$3389 "Straight Waveguide" sch_x=-27 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1696 N$3392 N$3391 "Straight Waveguide" sch_x=-27 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1697 N$3394 N$3393 "Straight Waveguide" sch_x=-27 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1698 N$3396 N$3395 "Straight Waveguide" sch_x=-27 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1699 N$3398 N$3397 "Straight Waveguide" sch_x=-27 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1700 N$3400 N$3399 "Straight Waveguide" sch_x=-27 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1701 N$3402 N$3401 "Straight Waveguide" sch_x=-27 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1702 N$3404 N$3403 "Straight Waveguide" sch_x=-27 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1703 N$3406 N$3405 "Straight Waveguide" sch_x=-27 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1704 N$3408 N$3407 "Straight Waveguide" sch_x=-27 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1705 N$3410 N$3409 "Straight Waveguide" sch_x=-27 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1706 N$3412 N$3411 "Straight Waveguide" sch_x=-27 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1707 N$3414 N$3413 "Straight Waveguide" sch_x=-25 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1708 N$3416 N$3415 "Straight Waveguide" sch_x=-25 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1709 N$3418 N$3417 "Straight Waveguide" sch_x=-25 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1710 N$3420 N$3419 "Straight Waveguide" sch_x=-25 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1711 N$3422 N$3421 "Straight Waveguide" sch_x=-25 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1712 N$3424 N$3423 "Straight Waveguide" sch_x=-25 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1713 N$3426 N$3425 "Straight Waveguide" sch_x=-25 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1714 N$3428 N$3427 "Straight Waveguide" sch_x=-25 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1715 N$3430 N$3429 "Straight Waveguide" sch_x=-25 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1716 N$3432 N$3431 "Straight Waveguide" sch_x=-25 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1717 N$3434 N$3433 "Straight Waveguide" sch_x=-23 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1718 N$3436 N$3435 "Straight Waveguide" sch_x=-23 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1719 N$3438 N$3437 "Straight Waveguide" sch_x=-23 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1720 N$3440 N$3439 "Straight Waveguide" sch_x=-23 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1721 N$3442 N$3441 "Straight Waveguide" sch_x=-23 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1722 N$3444 N$3443 "Straight Waveguide" sch_x=-23 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1723 N$3446 N$3445 "Straight Waveguide" sch_x=-23 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1724 N$3448 N$3447 "Straight Waveguide" sch_x=-23 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1725 N$3450 N$3449 "Straight Waveguide" sch_x=-21 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1726 N$3452 N$3451 "Straight Waveguide" sch_x=-21 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1727 N$3454 N$3453 "Straight Waveguide" sch_x=-21 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1728 N$3456 N$3455 "Straight Waveguide" sch_x=-21 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1729 N$3458 N$3457 "Straight Waveguide" sch_x=-21 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1730 N$3460 N$3459 "Straight Waveguide" sch_x=-21 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1731 N$3462 N$3461 "Straight Waveguide" sch_x=-19 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1732 N$3464 N$3463 "Straight Waveguide" sch_x=-19 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1733 N$3466 N$3465 "Straight Waveguide" sch_x=-19 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1734 N$3468 N$3467 "Straight Waveguide" sch_x=-19 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1735 N$3470 N$3469 "Straight Waveguide" sch_x=-17 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1736 N$3472 N$3471 "Straight Waveguide" sch_x=-17 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1737 N$3473 N$3474 "Straight Waveguide" sch_x=-21 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1738 N$3475 N$3476 "Straight Waveguide" sch_x=-20 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1739 N$3477 N$3478 "Straight Waveguide" sch_x=-19 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1740 N$3479 N$3480 "Straight Waveguide" sch_x=-18 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1741 N$3481 N$3482 "Straight Waveguide" sch_x=-17 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1742 N$3483 N$3484 "Straight Waveguide" sch_x=-16 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1743 N$3485 N$3486 "Straight Waveguide" sch_x=-15 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1744 N$3487 N$3488 "Straight Waveguide" sch_x=-15 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1745 N$3489 N$3490 "Straight Waveguide" sch_x=-16 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1746 N$3491 N$3492 "Straight Waveguide" sch_x=-17 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1747 N$3493 N$3494 "Straight Waveguide" sch_x=-18 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1748 N$3495 N$3496 "Straight Waveguide" sch_x=-19 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1749 N$3497 N$3498 "Straight Waveguide" sch_x=-20 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1750 N$3499 N$3500 "Straight Waveguide" sch_x=-21 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1751 N$3501 N$3502 "Straight Waveguide" sch_x=-22 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1752 N$3503 N$3504 "Straight Waveguide" sch_x=-22 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1753 N$3505 N$3506 "Straight Waveguide" sch_x=29 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1754 N$3507 N$3508 "Straight Waveguide" sch_x=29 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1755 N$3509 N$3510 "Straight Waveguide" sch_x=29 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1756 N$3511 N$3512 "Straight Waveguide" sch_x=29 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1757 N$3513 N$3514 "Straight Waveguide" sch_x=29 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1758 N$3515 N$3516 "Straight Waveguide" sch_x=29 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1759 N$3517 N$3518 "Straight Waveguide" sch_x=29 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1760 N$3519 N$3520 "Straight Waveguide" sch_x=29 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1761 N$3521 N$3522 "Straight Waveguide" sch_x=29 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1762 N$3523 N$3524 "Straight Waveguide" sch_x=29 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1763 N$3525 N$3526 "Straight Waveguide" sch_x=29 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1764 N$3527 N$3528 "Straight Waveguide" sch_x=29 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1765 N$3529 N$3530 "Straight Waveguide" sch_x=29 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1766 N$3531 N$3532 "Straight Waveguide" sch_x=29 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1767 N$3533 N$3534 "Straight Waveguide" sch_x=27 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1768 N$3535 N$3536 "Straight Waveguide" sch_x=27 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1769 N$3537 N$3538 "Straight Waveguide" sch_x=27 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1770 N$3539 N$3540 "Straight Waveguide" sch_x=27 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1771 N$3541 N$3542 "Straight Waveguide" sch_x=27 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1772 N$3543 N$3544 "Straight Waveguide" sch_x=27 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1773 N$3545 N$3546 "Straight Waveguide" sch_x=27 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1774 N$3547 N$3548 "Straight Waveguide" sch_x=27 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1775 N$3549 N$3550 "Straight Waveguide" sch_x=27 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1776 N$3551 N$3552 "Straight Waveguide" sch_x=27 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1777 N$3553 N$3554 "Straight Waveguide" sch_x=27 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1778 N$3555 N$3556 "Straight Waveguide" sch_x=27 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1779 N$3557 N$3558 "Straight Waveguide" sch_x=25 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1780 N$3559 N$3560 "Straight Waveguide" sch_x=25 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1781 N$3561 N$3562 "Straight Waveguide" sch_x=25 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1782 N$3563 N$3564 "Straight Waveguide" sch_x=25 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1783 N$3565 N$3566 "Straight Waveguide" sch_x=25 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1784 N$3567 N$3568 "Straight Waveguide" sch_x=25 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1785 N$3569 N$3570 "Straight Waveguide" sch_x=25 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1786 N$3571 N$3572 "Straight Waveguide" sch_x=25 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1787 N$3573 N$3574 "Straight Waveguide" sch_x=25 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1788 N$3575 N$3576 "Straight Waveguide" sch_x=25 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1789 N$3577 N$3578 "Straight Waveguide" sch_x=23 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1790 N$3579 N$3580 "Straight Waveguide" sch_x=23 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1791 N$3581 N$3582 "Straight Waveguide" sch_x=23 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1792 N$3583 N$3584 "Straight Waveguide" sch_x=23 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1793 N$3585 N$3586 "Straight Waveguide" sch_x=23 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1794 N$3587 N$3588 "Straight Waveguide" sch_x=23 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1795 N$3589 N$3590 "Straight Waveguide" sch_x=23 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1796 N$3591 N$3592 "Straight Waveguide" sch_x=23 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1797 N$3593 N$3594 "Straight Waveguide" sch_x=21 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1798 N$3595 N$3596 "Straight Waveguide" sch_x=21 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1799 N$3597 N$3598 "Straight Waveguide" sch_x=21 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1800 N$3599 N$3600 "Straight Waveguide" sch_x=21 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1801 N$3601 N$3602 "Straight Waveguide" sch_x=21 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1802 N$3603 N$3604 "Straight Waveguide" sch_x=21 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1803 N$3605 N$3606 "Straight Waveguide" sch_x=19 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1804 N$3607 N$3608 "Straight Waveguide" sch_x=19 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1805 N$3609 N$3610 "Straight Waveguide" sch_x=19 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1806 N$3611 N$3612 "Straight Waveguide" sch_x=19 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1807 N$3613 N$3614 "Straight Waveguide" sch_x=17 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1808 N$3615 N$3616 "Straight Waveguide" sch_x=17 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1809 N$3618 N$3617 "Straight Waveguide" sch_x=21 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1810 N$3620 N$3619 "Straight Waveguide" sch_x=20 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1811 N$3622 N$3621 "Straight Waveguide" sch_x=19 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1812 N$3624 N$3623 "Straight Waveguide" sch_x=18 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1813 N$3626 N$3625 "Straight Waveguide" sch_x=17 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1814 N$3628 N$3627 "Straight Waveguide" sch_x=16 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1815 N$3630 N$3629 "Straight Waveguide" sch_x=15 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1816 N$3632 N$3631 "Straight Waveguide" sch_x=15 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1817 N$3634 N$3633 "Straight Waveguide" sch_x=16 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1818 N$3636 N$3635 "Straight Waveguide" sch_x=17 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1819 N$3638 N$3637 "Straight Waveguide" sch_x=18 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1820 N$3640 N$3639 "Straight Waveguide" sch_x=19 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1821 N$3642 N$3641 "Straight Waveguide" sch_x=20 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1822 N$3644 N$3643 "Straight Waveguide" sch_x=21 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1823 N$3646 N$3645 "Straight Waveguide" sch_x=22 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1824 N$3648 N$3647 "Straight Waveguide" sch_x=22 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1825 N$3650 N$3649 "Straight Waveguide" sch_x=-61 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1826 N$3652 N$3651 "Straight Waveguide" sch_x=-61 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1827 N$3654 N$3653 "Straight Waveguide" sch_x=-61 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1828 N$3656 N$3655 "Straight Waveguide" sch_x=-61 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1829 N$3658 N$3657 "Straight Waveguide" sch_x=-61 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1830 N$3660 N$3659 "Straight Waveguide" sch_x=-61 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1831 N$3662 N$3661 "Straight Waveguide" sch_x=-61 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1832 N$3664 N$3663 "Straight Waveguide" sch_x=-61 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1833 N$3666 N$3665 "Straight Waveguide" sch_x=-61 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1834 N$3668 N$3667 "Straight Waveguide" sch_x=-61 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1835 N$3670 N$3669 "Straight Waveguide" sch_x=-61 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1836 N$3672 N$3671 "Straight Waveguide" sch_x=-61 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1837 N$3674 N$3673 "Straight Waveguide" sch_x=-61 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1838 N$3676 N$3675 "Straight Waveguide" sch_x=-61 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1839 N$3678 N$3677 "Straight Waveguide" sch_x=-61 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1840 N$3680 N$3679 "Straight Waveguide" sch_x=-61 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1841 N$3682 N$3681 "Straight Waveguide" sch_x=-61 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1842 N$3684 N$3683 "Straight Waveguide" sch_x=-61 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1843 N$3686 N$3685 "Straight Waveguide" sch_x=-61 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1844 N$3688 N$3687 "Straight Waveguide" sch_x=-61 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1845 N$3690 N$3689 "Straight Waveguide" sch_x=-61 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1846 N$3692 N$3691 "Straight Waveguide" sch_x=-61 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1847 N$3694 N$3693 "Straight Waveguide" sch_x=-61 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1848 N$3696 N$3695 "Straight Waveguide" sch_x=-61 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1849 N$3698 N$3697 "Straight Waveguide" sch_x=-61 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1850 N$3700 N$3699 "Straight Waveguide" sch_x=-61 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1851 N$3702 N$3701 "Straight Waveguide" sch_x=-61 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1852 N$3704 N$3703 "Straight Waveguide" sch_x=-61 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1853 N$3706 N$3705 "Straight Waveguide" sch_x=-61 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1854 N$3708 N$3707 "Straight Waveguide" sch_x=-61 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1855 N$3710 N$3709 "Straight Waveguide" sch_x=-59 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1856 N$3712 N$3711 "Straight Waveguide" sch_x=-59 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1857 N$3714 N$3713 "Straight Waveguide" sch_x=-59 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1858 N$3716 N$3715 "Straight Waveguide" sch_x=-59 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1859 N$3718 N$3717 "Straight Waveguide" sch_x=-59 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1860 N$3720 N$3719 "Straight Waveguide" sch_x=-59 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1861 N$3722 N$3721 "Straight Waveguide" sch_x=-59 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1862 N$3724 N$3723 "Straight Waveguide" sch_x=-59 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1863 N$3726 N$3725 "Straight Waveguide" sch_x=-59 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1864 N$3728 N$3727 "Straight Waveguide" sch_x=-59 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1865 N$3730 N$3729 "Straight Waveguide" sch_x=-59 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1866 N$3732 N$3731 "Straight Waveguide" sch_x=-59 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1867 N$3734 N$3733 "Straight Waveguide" sch_x=-59 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1868 N$3736 N$3735 "Straight Waveguide" sch_x=-59 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1869 N$3738 N$3737 "Straight Waveguide" sch_x=-59 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1870 N$3740 N$3739 "Straight Waveguide" sch_x=-59 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1871 N$3742 N$3741 "Straight Waveguide" sch_x=-59 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1872 N$3744 N$3743 "Straight Waveguide" sch_x=-59 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1873 N$3746 N$3745 "Straight Waveguide" sch_x=-59 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1874 N$3748 N$3747 "Straight Waveguide" sch_x=-59 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1875 N$3750 N$3749 "Straight Waveguide" sch_x=-59 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1876 N$3752 N$3751 "Straight Waveguide" sch_x=-59 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1877 N$3754 N$3753 "Straight Waveguide" sch_x=-59 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1878 N$3756 N$3755 "Straight Waveguide" sch_x=-59 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1879 N$3758 N$3757 "Straight Waveguide" sch_x=-59 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1880 N$3760 N$3759 "Straight Waveguide" sch_x=-59 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1881 N$3762 N$3761 "Straight Waveguide" sch_x=-59 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1882 N$3764 N$3763 "Straight Waveguide" sch_x=-59 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1883 N$3766 N$3765 "Straight Waveguide" sch_x=-57 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1884 N$3768 N$3767 "Straight Waveguide" sch_x=-57 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1885 N$3770 N$3769 "Straight Waveguide" sch_x=-57 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1886 N$3772 N$3771 "Straight Waveguide" sch_x=-57 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1887 N$3774 N$3773 "Straight Waveguide" sch_x=-57 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1888 N$3776 N$3775 "Straight Waveguide" sch_x=-57 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1889 N$3778 N$3777 "Straight Waveguide" sch_x=-57 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1890 N$3780 N$3779 "Straight Waveguide" sch_x=-57 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1891 N$3782 N$3781 "Straight Waveguide" sch_x=-57 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1892 N$3784 N$3783 "Straight Waveguide" sch_x=-57 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1893 N$3786 N$3785 "Straight Waveguide" sch_x=-57 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1894 N$3788 N$3787 "Straight Waveguide" sch_x=-57 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1895 N$3790 N$3789 "Straight Waveguide" sch_x=-57 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1896 N$3792 N$3791 "Straight Waveguide" sch_x=-57 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1897 N$3794 N$3793 "Straight Waveguide" sch_x=-57 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1898 N$3796 N$3795 "Straight Waveguide" sch_x=-57 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1899 N$3798 N$3797 "Straight Waveguide" sch_x=-57 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1900 N$3800 N$3799 "Straight Waveguide" sch_x=-57 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1901 N$3802 N$3801 "Straight Waveguide" sch_x=-57 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1902 N$3804 N$3803 "Straight Waveguide" sch_x=-57 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1903 N$3806 N$3805 "Straight Waveguide" sch_x=-57 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1904 N$3808 N$3807 "Straight Waveguide" sch_x=-57 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1905 N$3810 N$3809 "Straight Waveguide" sch_x=-57 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1906 N$3812 N$3811 "Straight Waveguide" sch_x=-57 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1907 N$3814 N$3813 "Straight Waveguide" sch_x=-57 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1908 N$3816 N$3815 "Straight Waveguide" sch_x=-57 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1909 N$3818 N$3817 "Straight Waveguide" sch_x=-55 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1910 N$3820 N$3819 "Straight Waveguide" sch_x=-55 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1911 N$3822 N$3821 "Straight Waveguide" sch_x=-55 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1912 N$3824 N$3823 "Straight Waveguide" sch_x=-55 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1913 N$3826 N$3825 "Straight Waveguide" sch_x=-55 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1914 N$3828 N$3827 "Straight Waveguide" sch_x=-55 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1915 N$3830 N$3829 "Straight Waveguide" sch_x=-55 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1916 N$3832 N$3831 "Straight Waveguide" sch_x=-55 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1917 N$3834 N$3833 "Straight Waveguide" sch_x=-55 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1918 N$3836 N$3835 "Straight Waveguide" sch_x=-55 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1919 N$3838 N$3837 "Straight Waveguide" sch_x=-55 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1920 N$3840 N$3839 "Straight Waveguide" sch_x=-55 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1921 N$3842 N$3841 "Straight Waveguide" sch_x=-55 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1922 N$3844 N$3843 "Straight Waveguide" sch_x=-55 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1923 N$3846 N$3845 "Straight Waveguide" sch_x=-55 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1924 N$3848 N$3847 "Straight Waveguide" sch_x=-55 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1925 N$3850 N$3849 "Straight Waveguide" sch_x=-55 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1926 N$3852 N$3851 "Straight Waveguide" sch_x=-55 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1927 N$3854 N$3853 "Straight Waveguide" sch_x=-55 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1928 N$3856 N$3855 "Straight Waveguide" sch_x=-55 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1929 N$3858 N$3857 "Straight Waveguide" sch_x=-55 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1930 N$3860 N$3859 "Straight Waveguide" sch_x=-55 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1931 N$3862 N$3861 "Straight Waveguide" sch_x=-55 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1932 N$3864 N$3863 "Straight Waveguide" sch_x=-55 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1933 N$3866 N$3865 "Straight Waveguide" sch_x=-53 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1934 N$3868 N$3867 "Straight Waveguide" sch_x=-53 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1935 N$3870 N$3869 "Straight Waveguide" sch_x=-53 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1936 N$3872 N$3871 "Straight Waveguide" sch_x=-53 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1937 N$3874 N$3873 "Straight Waveguide" sch_x=-53 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1938 N$3876 N$3875 "Straight Waveguide" sch_x=-53 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1939 N$3878 N$3877 "Straight Waveguide" sch_x=-53 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1940 N$3880 N$3879 "Straight Waveguide" sch_x=-53 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1941 N$3882 N$3881 "Straight Waveguide" sch_x=-53 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1942 N$3884 N$3883 "Straight Waveguide" sch_x=-53 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1943 N$3886 N$3885 "Straight Waveguide" sch_x=-53 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1944 N$3888 N$3887 "Straight Waveguide" sch_x=-53 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1945 N$3890 N$3889 "Straight Waveguide" sch_x=-53 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1946 N$3892 N$3891 "Straight Waveguide" sch_x=-53 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1947 N$3894 N$3893 "Straight Waveguide" sch_x=-53 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1948 N$3896 N$3895 "Straight Waveguide" sch_x=-53 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1949 N$3898 N$3897 "Straight Waveguide" sch_x=-53 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1950 N$3900 N$3899 "Straight Waveguide" sch_x=-53 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1951 N$3902 N$3901 "Straight Waveguide" sch_x=-53 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1952 N$3904 N$3903 "Straight Waveguide" sch_x=-53 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1953 N$3906 N$3905 "Straight Waveguide" sch_x=-53 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1954 N$3908 N$3907 "Straight Waveguide" sch_x=-53 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1955 N$3910 N$3909 "Straight Waveguide" sch_x=-51 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1956 N$3912 N$3911 "Straight Waveguide" sch_x=-51 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1957 N$3914 N$3913 "Straight Waveguide" sch_x=-51 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1958 N$3916 N$3915 "Straight Waveguide" sch_x=-51 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1959 N$3918 N$3917 "Straight Waveguide" sch_x=-51 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1960 N$3920 N$3919 "Straight Waveguide" sch_x=-51 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1961 N$3922 N$3921 "Straight Waveguide" sch_x=-51 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1962 N$3924 N$3923 "Straight Waveguide" sch_x=-51 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1963 N$3926 N$3925 "Straight Waveguide" sch_x=-51 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1964 N$3928 N$3927 "Straight Waveguide" sch_x=-51 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1965 N$3930 N$3929 "Straight Waveguide" sch_x=-51 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1966 N$3932 N$3931 "Straight Waveguide" sch_x=-51 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1967 N$3934 N$3933 "Straight Waveguide" sch_x=-51 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1968 N$3936 N$3935 "Straight Waveguide" sch_x=-51 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1969 N$3938 N$3937 "Straight Waveguide" sch_x=-51 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1970 N$3940 N$3939 "Straight Waveguide" sch_x=-51 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1971 N$3942 N$3941 "Straight Waveguide" sch_x=-51 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1972 N$3944 N$3943 "Straight Waveguide" sch_x=-51 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1973 N$3946 N$3945 "Straight Waveguide" sch_x=-51 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1974 N$3948 N$3947 "Straight Waveguide" sch_x=-51 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1975 N$3950 N$3949 "Straight Waveguide" sch_x=-49 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1976 N$3952 N$3951 "Straight Waveguide" sch_x=-49 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1977 N$3954 N$3953 "Straight Waveguide" sch_x=-49 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1978 N$3956 N$3955 "Straight Waveguide" sch_x=-49 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1979 N$3958 N$3957 "Straight Waveguide" sch_x=-49 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1980 N$3960 N$3959 "Straight Waveguide" sch_x=-49 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1981 N$3962 N$3961 "Straight Waveguide" sch_x=-49 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1982 N$3964 N$3963 "Straight Waveguide" sch_x=-49 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1983 N$3966 N$3965 "Straight Waveguide" sch_x=-49 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1984 N$3968 N$3967 "Straight Waveguide" sch_x=-49 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1985 N$3970 N$3969 "Straight Waveguide" sch_x=-49 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1986 N$3972 N$3971 "Straight Waveguide" sch_x=-49 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1987 N$3974 N$3973 "Straight Waveguide" sch_x=-49 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1988 N$3976 N$3975 "Straight Waveguide" sch_x=-49 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1989 N$3978 N$3977 "Straight Waveguide" sch_x=-49 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1990 N$3980 N$3979 "Straight Waveguide" sch_x=-49 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1991 N$3982 N$3981 "Straight Waveguide" sch_x=-49 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1992 N$3984 N$3983 "Straight Waveguide" sch_x=-49 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1993 N$3986 N$3985 "Straight Waveguide" sch_x=-47 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1994 N$3988 N$3987 "Straight Waveguide" sch_x=-47 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1995 N$3990 N$3989 "Straight Waveguide" sch_x=-47 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1996 N$3992 N$3991 "Straight Waveguide" sch_x=-47 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1997 N$3994 N$3993 "Straight Waveguide" sch_x=-47 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1998 N$3996 N$3995 "Straight Waveguide" sch_x=-47 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W1999 N$3998 N$3997 "Straight Waveguide" sch_x=-47 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2000 N$4000 N$3999 "Straight Waveguide" sch_x=-47 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2001 N$4002 N$4001 "Straight Waveguide" sch_x=-47 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2002 N$4004 N$4003 "Straight Waveguide" sch_x=-47 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2003 N$4006 N$4005 "Straight Waveguide" sch_x=-47 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2004 N$4008 N$4007 "Straight Waveguide" sch_x=-47 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2005 N$4010 N$4009 "Straight Waveguide" sch_x=-47 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2006 N$4012 N$4011 "Straight Waveguide" sch_x=-47 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2007 N$4014 N$4013 "Straight Waveguide" sch_x=-47 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2008 N$4016 N$4015 "Straight Waveguide" sch_x=-47 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2009 N$4018 N$4017 "Straight Waveguide" sch_x=-45 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2010 N$4020 N$4019 "Straight Waveguide" sch_x=-45 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2011 N$4022 N$4021 "Straight Waveguide" sch_x=-45 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2012 N$4024 N$4023 "Straight Waveguide" sch_x=-45 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2013 N$4026 N$4025 "Straight Waveguide" sch_x=-45 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2014 N$4028 N$4027 "Straight Waveguide" sch_x=-45 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2015 N$4030 N$4029 "Straight Waveguide" sch_x=-45 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2016 N$4032 N$4031 "Straight Waveguide" sch_x=-45 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2017 N$4034 N$4033 "Straight Waveguide" sch_x=-45 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2018 N$4036 N$4035 "Straight Waveguide" sch_x=-45 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2019 N$4038 N$4037 "Straight Waveguide" sch_x=-45 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2020 N$4040 N$4039 "Straight Waveguide" sch_x=-45 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2021 N$4042 N$4041 "Straight Waveguide" sch_x=-45 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2022 N$4044 N$4043 "Straight Waveguide" sch_x=-45 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2023 N$4046 N$4045 "Straight Waveguide" sch_x=-43 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2024 N$4048 N$4047 "Straight Waveguide" sch_x=-43 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2025 N$4050 N$4049 "Straight Waveguide" sch_x=-43 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2026 N$4052 N$4051 "Straight Waveguide" sch_x=-43 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2027 N$4054 N$4053 "Straight Waveguide" sch_x=-43 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2028 N$4056 N$4055 "Straight Waveguide" sch_x=-43 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2029 N$4058 N$4057 "Straight Waveguide" sch_x=-43 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2030 N$4060 N$4059 "Straight Waveguide" sch_x=-43 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2031 N$4062 N$4061 "Straight Waveguide" sch_x=-43 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2032 N$4064 N$4063 "Straight Waveguide" sch_x=-43 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2033 N$4066 N$4065 "Straight Waveguide" sch_x=-43 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2034 N$4068 N$4067 "Straight Waveguide" sch_x=-43 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2035 N$4070 N$4069 "Straight Waveguide" sch_x=-41 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2036 N$4072 N$4071 "Straight Waveguide" sch_x=-41 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2037 N$4074 N$4073 "Straight Waveguide" sch_x=-41 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2038 N$4076 N$4075 "Straight Waveguide" sch_x=-41 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2039 N$4078 N$4077 "Straight Waveguide" sch_x=-41 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2040 N$4080 N$4079 "Straight Waveguide" sch_x=-41 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2041 N$4082 N$4081 "Straight Waveguide" sch_x=-41 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2042 N$4084 N$4083 "Straight Waveguide" sch_x=-41 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2043 N$4086 N$4085 "Straight Waveguide" sch_x=-41 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2044 N$4088 N$4087 "Straight Waveguide" sch_x=-41 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2045 N$4090 N$4089 "Straight Waveguide" sch_x=-39 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2046 N$4092 N$4091 "Straight Waveguide" sch_x=-39 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2047 N$4094 N$4093 "Straight Waveguide" sch_x=-39 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2048 N$4096 N$4095 "Straight Waveguide" sch_x=-39 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2049 N$4098 N$4097 "Straight Waveguide" sch_x=-39 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2050 N$4100 N$4099 "Straight Waveguide" sch_x=-39 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2051 N$4102 N$4101 "Straight Waveguide" sch_x=-39 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2052 N$4104 N$4103 "Straight Waveguide" sch_x=-39 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2053 N$4106 N$4105 "Straight Waveguide" sch_x=-37 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2054 N$4108 N$4107 "Straight Waveguide" sch_x=-37 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2055 N$4110 N$4109 "Straight Waveguide" sch_x=-37 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2056 N$4112 N$4111 "Straight Waveguide" sch_x=-37 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2057 N$4114 N$4113 "Straight Waveguide" sch_x=-37 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2058 N$4116 N$4115 "Straight Waveguide" sch_x=-37 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2059 N$4118 N$4117 "Straight Waveguide" sch_x=-35 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2060 N$4120 N$4119 "Straight Waveguide" sch_x=-35 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2061 N$4122 N$4121 "Straight Waveguide" sch_x=-35 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2062 N$4124 N$4123 "Straight Waveguide" sch_x=-35 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2063 N$4126 N$4125 "Straight Waveguide" sch_x=-33 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2064 N$4128 N$4127 "Straight Waveguide" sch_x=-33 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2065 N$4129 N$4130 "Straight Waveguide" sch_x=-45 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2066 N$4131 N$4132 "Straight Waveguide" sch_x=-44 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2067 N$4133 N$4134 "Straight Waveguide" sch_x=-43 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2068 N$4135 N$4136 "Straight Waveguide" sch_x=-42 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2069 N$4137 N$4138 "Straight Waveguide" sch_x=-41 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2070 N$4139 N$4140 "Straight Waveguide" sch_x=-40 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2071 N$4141 N$4142 "Straight Waveguide" sch_x=-39 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2072 N$4143 N$4144 "Straight Waveguide" sch_x=-38 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2073 N$4145 N$4146 "Straight Waveguide" sch_x=-37 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2074 N$4147 N$4148 "Straight Waveguide" sch_x=-36 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2075 N$4149 N$4150 "Straight Waveguide" sch_x=-35 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2076 N$4151 N$4152 "Straight Waveguide" sch_x=-34 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2077 N$4153 N$4154 "Straight Waveguide" sch_x=-33 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2078 N$4155 N$4156 "Straight Waveguide" sch_x=-32 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2079 N$4157 N$4158 "Straight Waveguide" sch_x=-31 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2080 N$4159 N$4160 "Straight Waveguide" sch_x=-31 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2081 N$4161 N$4162 "Straight Waveguide" sch_x=-32 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2082 N$4163 N$4164 "Straight Waveguide" sch_x=-33 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2083 N$4165 N$4166 "Straight Waveguide" sch_x=-34 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2084 N$4167 N$4168 "Straight Waveguide" sch_x=-35 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2085 N$4169 N$4170 "Straight Waveguide" sch_x=-36 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2086 N$4171 N$4172 "Straight Waveguide" sch_x=-37 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2087 N$4173 N$4174 "Straight Waveguide" sch_x=-38 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2088 N$4175 N$4176 "Straight Waveguide" sch_x=-39 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2089 N$4177 N$4178 "Straight Waveguide" sch_x=-40 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2090 N$4179 N$4180 "Straight Waveguide" sch_x=-41 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2091 N$4181 N$4182 "Straight Waveguide" sch_x=-42 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2092 N$4183 N$4184 "Straight Waveguide" sch_x=-43 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2093 N$4185 N$4186 "Straight Waveguide" sch_x=-44 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2094 N$4187 N$4188 "Straight Waveguide" sch_x=-45 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2095 N$4189 N$4190 "Straight Waveguide" sch_x=-46 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2096 N$4191 N$4192 "Straight Waveguide" sch_x=-46 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2097 N$4193 N$4194 "Straight Waveguide" sch_x=61 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2098 N$4195 N$4196 "Straight Waveguide" sch_x=61 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2099 N$4197 N$4198 "Straight Waveguide" sch_x=61 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2100 N$4199 N$4200 "Straight Waveguide" sch_x=61 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2101 N$4201 N$4202 "Straight Waveguide" sch_x=61 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2102 N$4203 N$4204 "Straight Waveguide" sch_x=61 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2103 N$4205 N$4206 "Straight Waveguide" sch_x=61 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2104 N$4207 N$4208 "Straight Waveguide" sch_x=61 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2105 N$4209 N$4210 "Straight Waveguide" sch_x=61 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2106 N$4211 N$4212 "Straight Waveguide" sch_x=61 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2107 N$4213 N$4214 "Straight Waveguide" sch_x=61 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2108 N$4215 N$4216 "Straight Waveguide" sch_x=61 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2109 N$4217 N$4218 "Straight Waveguide" sch_x=61 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2110 N$4219 N$4220 "Straight Waveguide" sch_x=61 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2111 N$4221 N$4222 "Straight Waveguide" sch_x=61 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2112 N$4223 N$4224 "Straight Waveguide" sch_x=61 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2113 N$4225 N$4226 "Straight Waveguide" sch_x=61 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2114 N$4227 N$4228 "Straight Waveguide" sch_x=61 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2115 N$4229 N$4230 "Straight Waveguide" sch_x=61 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2116 N$4231 N$4232 "Straight Waveguide" sch_x=61 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2117 N$4233 N$4234 "Straight Waveguide" sch_x=61 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2118 N$4235 N$4236 "Straight Waveguide" sch_x=61 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2119 N$4237 N$4238 "Straight Waveguide" sch_x=61 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2120 N$4239 N$4240 "Straight Waveguide" sch_x=61 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2121 N$4241 N$4242 "Straight Waveguide" sch_x=61 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2122 N$4243 N$4244 "Straight Waveguide" sch_x=61 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2123 N$4245 N$4246 "Straight Waveguide" sch_x=61 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2124 N$4247 N$4248 "Straight Waveguide" sch_x=61 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2125 N$4249 N$4250 "Straight Waveguide" sch_x=61 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2126 N$4251 N$4252 "Straight Waveguide" sch_x=61 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2127 N$4253 N$4254 "Straight Waveguide" sch_x=59 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2128 N$4255 N$4256 "Straight Waveguide" sch_x=59 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2129 N$4257 N$4258 "Straight Waveguide" sch_x=59 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2130 N$4259 N$4260 "Straight Waveguide" sch_x=59 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2131 N$4261 N$4262 "Straight Waveguide" sch_x=59 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2132 N$4263 N$4264 "Straight Waveguide" sch_x=59 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2133 N$4265 N$4266 "Straight Waveguide" sch_x=59 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2134 N$4267 N$4268 "Straight Waveguide" sch_x=59 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2135 N$4269 N$4270 "Straight Waveguide" sch_x=59 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2136 N$4271 N$4272 "Straight Waveguide" sch_x=59 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2137 N$4273 N$4274 "Straight Waveguide" sch_x=59 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2138 N$4275 N$4276 "Straight Waveguide" sch_x=59 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2139 N$4277 N$4278 "Straight Waveguide" sch_x=59 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2140 N$4279 N$4280 "Straight Waveguide" sch_x=59 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2141 N$4281 N$4282 "Straight Waveguide" sch_x=59 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2142 N$4283 N$4284 "Straight Waveguide" sch_x=59 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2143 N$4285 N$4286 "Straight Waveguide" sch_x=59 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2144 N$4287 N$4288 "Straight Waveguide" sch_x=59 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2145 N$4289 N$4290 "Straight Waveguide" sch_x=59 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2146 N$4291 N$4292 "Straight Waveguide" sch_x=59 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2147 N$4293 N$4294 "Straight Waveguide" sch_x=59 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2148 N$4295 N$4296 "Straight Waveguide" sch_x=59 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2149 N$4297 N$4298 "Straight Waveguide" sch_x=59 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2150 N$4299 N$4300 "Straight Waveguide" sch_x=59 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2151 N$4301 N$4302 "Straight Waveguide" sch_x=59 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2152 N$4303 N$4304 "Straight Waveguide" sch_x=59 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2153 N$4305 N$4306 "Straight Waveguide" sch_x=59 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2154 N$4307 N$4308 "Straight Waveguide" sch_x=59 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2155 N$4309 N$4310 "Straight Waveguide" sch_x=57 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2156 N$4311 N$4312 "Straight Waveguide" sch_x=57 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2157 N$4313 N$4314 "Straight Waveguide" sch_x=57 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2158 N$4315 N$4316 "Straight Waveguide" sch_x=57 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2159 N$4317 N$4318 "Straight Waveguide" sch_x=57 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2160 N$4319 N$4320 "Straight Waveguide" sch_x=57 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2161 N$4321 N$4322 "Straight Waveguide" sch_x=57 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2162 N$4323 N$4324 "Straight Waveguide" sch_x=57 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2163 N$4325 N$4326 "Straight Waveguide" sch_x=57 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2164 N$4327 N$4328 "Straight Waveguide" sch_x=57 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2165 N$4329 N$4330 "Straight Waveguide" sch_x=57 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2166 N$4331 N$4332 "Straight Waveguide" sch_x=57 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2167 N$4333 N$4334 "Straight Waveguide" sch_x=57 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2168 N$4335 N$4336 "Straight Waveguide" sch_x=57 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2169 N$4337 N$4338 "Straight Waveguide" sch_x=57 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2170 N$4339 N$4340 "Straight Waveguide" sch_x=57 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2171 N$4341 N$4342 "Straight Waveguide" sch_x=57 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2172 N$4343 N$4344 "Straight Waveguide" sch_x=57 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2173 N$4345 N$4346 "Straight Waveguide" sch_x=57 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2174 N$4347 N$4348 "Straight Waveguide" sch_x=57 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2175 N$4349 N$4350 "Straight Waveguide" sch_x=57 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2176 N$4351 N$4352 "Straight Waveguide" sch_x=57 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2177 N$4353 N$4354 "Straight Waveguide" sch_x=57 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2178 N$4355 N$4356 "Straight Waveguide" sch_x=57 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2179 N$4357 N$4358 "Straight Waveguide" sch_x=57 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2180 N$4359 N$4360 "Straight Waveguide" sch_x=57 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2181 N$4361 N$4362 "Straight Waveguide" sch_x=55 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2182 N$4363 N$4364 "Straight Waveguide" sch_x=55 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2183 N$4365 N$4366 "Straight Waveguide" sch_x=55 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2184 N$4367 N$4368 "Straight Waveguide" sch_x=55 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2185 N$4369 N$4370 "Straight Waveguide" sch_x=55 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2186 N$4371 N$4372 "Straight Waveguide" sch_x=55 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2187 N$4373 N$4374 "Straight Waveguide" sch_x=55 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2188 N$4375 N$4376 "Straight Waveguide" sch_x=55 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2189 N$4377 N$4378 "Straight Waveguide" sch_x=55 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2190 N$4379 N$4380 "Straight Waveguide" sch_x=55 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2191 N$4381 N$4382 "Straight Waveguide" sch_x=55 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2192 N$4383 N$4384 "Straight Waveguide" sch_x=55 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2193 N$4385 N$4386 "Straight Waveguide" sch_x=55 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2194 N$4387 N$4388 "Straight Waveguide" sch_x=55 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2195 N$4389 N$4390 "Straight Waveguide" sch_x=55 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2196 N$4391 N$4392 "Straight Waveguide" sch_x=55 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2197 N$4393 N$4394 "Straight Waveguide" sch_x=55 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2198 N$4395 N$4396 "Straight Waveguide" sch_x=55 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2199 N$4397 N$4398 "Straight Waveguide" sch_x=55 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2200 N$4399 N$4400 "Straight Waveguide" sch_x=55 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2201 N$4401 N$4402 "Straight Waveguide" sch_x=55 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2202 N$4403 N$4404 "Straight Waveguide" sch_x=55 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2203 N$4405 N$4406 "Straight Waveguide" sch_x=55 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2204 N$4407 N$4408 "Straight Waveguide" sch_x=55 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2205 N$4409 N$4410 "Straight Waveguide" sch_x=53 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2206 N$4411 N$4412 "Straight Waveguide" sch_x=53 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2207 N$4413 N$4414 "Straight Waveguide" sch_x=53 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2208 N$4415 N$4416 "Straight Waveguide" sch_x=53 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2209 N$4417 N$4418 "Straight Waveguide" sch_x=53 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2210 N$4419 N$4420 "Straight Waveguide" sch_x=53 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2211 N$4421 N$4422 "Straight Waveguide" sch_x=53 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2212 N$4423 N$4424 "Straight Waveguide" sch_x=53 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2213 N$4425 N$4426 "Straight Waveguide" sch_x=53 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2214 N$4427 N$4428 "Straight Waveguide" sch_x=53 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2215 N$4429 N$4430 "Straight Waveguide" sch_x=53 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2216 N$4431 N$4432 "Straight Waveguide" sch_x=53 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2217 N$4433 N$4434 "Straight Waveguide" sch_x=53 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2218 N$4435 N$4436 "Straight Waveguide" sch_x=53 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2219 N$4437 N$4438 "Straight Waveguide" sch_x=53 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2220 N$4439 N$4440 "Straight Waveguide" sch_x=53 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2221 N$4441 N$4442 "Straight Waveguide" sch_x=53 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2222 N$4443 N$4444 "Straight Waveguide" sch_x=53 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2223 N$4445 N$4446 "Straight Waveguide" sch_x=53 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2224 N$4447 N$4448 "Straight Waveguide" sch_x=53 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2225 N$4449 N$4450 "Straight Waveguide" sch_x=53 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2226 N$4451 N$4452 "Straight Waveguide" sch_x=53 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2227 N$4453 N$4454 "Straight Waveguide" sch_x=51 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2228 N$4455 N$4456 "Straight Waveguide" sch_x=51 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2229 N$4457 N$4458 "Straight Waveguide" sch_x=51 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2230 N$4459 N$4460 "Straight Waveguide" sch_x=51 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2231 N$4461 N$4462 "Straight Waveguide" sch_x=51 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2232 N$4463 N$4464 "Straight Waveguide" sch_x=51 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2233 N$4465 N$4466 "Straight Waveguide" sch_x=51 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2234 N$4467 N$4468 "Straight Waveguide" sch_x=51 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2235 N$4469 N$4470 "Straight Waveguide" sch_x=51 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2236 N$4471 N$4472 "Straight Waveguide" sch_x=51 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2237 N$4473 N$4474 "Straight Waveguide" sch_x=51 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2238 N$4475 N$4476 "Straight Waveguide" sch_x=51 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2239 N$4477 N$4478 "Straight Waveguide" sch_x=51 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2240 N$4479 N$4480 "Straight Waveguide" sch_x=51 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2241 N$4481 N$4482 "Straight Waveguide" sch_x=51 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2242 N$4483 N$4484 "Straight Waveguide" sch_x=51 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2243 N$4485 N$4486 "Straight Waveguide" sch_x=51 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2244 N$4487 N$4488 "Straight Waveguide" sch_x=51 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2245 N$4489 N$4490 "Straight Waveguide" sch_x=51 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2246 N$4491 N$4492 "Straight Waveguide" sch_x=51 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2247 N$4493 N$4494 "Straight Waveguide" sch_x=49 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2248 N$4495 N$4496 "Straight Waveguide" sch_x=49 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2249 N$4497 N$4498 "Straight Waveguide" sch_x=49 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2250 N$4499 N$4500 "Straight Waveguide" sch_x=49 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2251 N$4501 N$4502 "Straight Waveguide" sch_x=49 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2252 N$4503 N$4504 "Straight Waveguide" sch_x=49 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2253 N$4505 N$4506 "Straight Waveguide" sch_x=49 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2254 N$4507 N$4508 "Straight Waveguide" sch_x=49 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2255 N$4509 N$4510 "Straight Waveguide" sch_x=49 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2256 N$4511 N$4512 "Straight Waveguide" sch_x=49 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2257 N$4513 N$4514 "Straight Waveguide" sch_x=49 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2258 N$4515 N$4516 "Straight Waveguide" sch_x=49 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2259 N$4517 N$4518 "Straight Waveguide" sch_x=49 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2260 N$4519 N$4520 "Straight Waveguide" sch_x=49 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2261 N$4521 N$4522 "Straight Waveguide" sch_x=49 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2262 N$4523 N$4524 "Straight Waveguide" sch_x=49 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2263 N$4525 N$4526 "Straight Waveguide" sch_x=49 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2264 N$4527 N$4528 "Straight Waveguide" sch_x=49 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2265 N$4529 N$4530 "Straight Waveguide" sch_x=47 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2266 N$4531 N$4532 "Straight Waveguide" sch_x=47 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2267 N$4533 N$4534 "Straight Waveguide" sch_x=47 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2268 N$4535 N$4536 "Straight Waveguide" sch_x=47 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2269 N$4537 N$4538 "Straight Waveguide" sch_x=47 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2270 N$4539 N$4540 "Straight Waveguide" sch_x=47 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2271 N$4541 N$4542 "Straight Waveguide" sch_x=47 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2272 N$4543 N$4544 "Straight Waveguide" sch_x=47 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2273 N$4545 N$4546 "Straight Waveguide" sch_x=47 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2274 N$4547 N$4548 "Straight Waveguide" sch_x=47 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2275 N$4549 N$4550 "Straight Waveguide" sch_x=47 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2276 N$4551 N$4552 "Straight Waveguide" sch_x=47 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2277 N$4553 N$4554 "Straight Waveguide" sch_x=47 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2278 N$4555 N$4556 "Straight Waveguide" sch_x=47 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2279 N$4557 N$4558 "Straight Waveguide" sch_x=47 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2280 N$4559 N$4560 "Straight Waveguide" sch_x=47 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2281 N$4561 N$4562 "Straight Waveguide" sch_x=45 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2282 N$4563 N$4564 "Straight Waveguide" sch_x=45 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2283 N$4565 N$4566 "Straight Waveguide" sch_x=45 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2284 N$4567 N$4568 "Straight Waveguide" sch_x=45 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2285 N$4569 N$4570 "Straight Waveguide" sch_x=45 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2286 N$4571 N$4572 "Straight Waveguide" sch_x=45 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2287 N$4573 N$4574 "Straight Waveguide" sch_x=45 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2288 N$4575 N$4576 "Straight Waveguide" sch_x=45 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2289 N$4577 N$4578 "Straight Waveguide" sch_x=45 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2290 N$4579 N$4580 "Straight Waveguide" sch_x=45 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2291 N$4581 N$4582 "Straight Waveguide" sch_x=45 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2292 N$4583 N$4584 "Straight Waveguide" sch_x=45 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2293 N$4585 N$4586 "Straight Waveguide" sch_x=45 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2294 N$4587 N$4588 "Straight Waveguide" sch_x=45 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2295 N$4589 N$4590 "Straight Waveguide" sch_x=43 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2296 N$4591 N$4592 "Straight Waveguide" sch_x=43 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2297 N$4593 N$4594 "Straight Waveguide" sch_x=43 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2298 N$4595 N$4596 "Straight Waveguide" sch_x=43 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2299 N$4597 N$4598 "Straight Waveguide" sch_x=43 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2300 N$4599 N$4600 "Straight Waveguide" sch_x=43 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2301 N$4601 N$4602 "Straight Waveguide" sch_x=43 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2302 N$4603 N$4604 "Straight Waveguide" sch_x=43 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2303 N$4605 N$4606 "Straight Waveguide" sch_x=43 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2304 N$4607 N$4608 "Straight Waveguide" sch_x=43 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2305 N$4609 N$4610 "Straight Waveguide" sch_x=43 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2306 N$4611 N$4612 "Straight Waveguide" sch_x=43 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2307 N$4613 N$4614 "Straight Waveguide" sch_x=41 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2308 N$4615 N$4616 "Straight Waveguide" sch_x=41 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2309 N$4617 N$4618 "Straight Waveguide" sch_x=41 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2310 N$4619 N$4620 "Straight Waveguide" sch_x=41 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2311 N$4621 N$4622 "Straight Waveguide" sch_x=41 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2312 N$4623 N$4624 "Straight Waveguide" sch_x=41 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2313 N$4625 N$4626 "Straight Waveguide" sch_x=41 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2314 N$4627 N$4628 "Straight Waveguide" sch_x=41 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2315 N$4629 N$4630 "Straight Waveguide" sch_x=41 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2316 N$4631 N$4632 "Straight Waveguide" sch_x=41 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2317 N$4633 N$4634 "Straight Waveguide" sch_x=39 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2318 N$4635 N$4636 "Straight Waveguide" sch_x=39 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2319 N$4637 N$4638 "Straight Waveguide" sch_x=39 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2320 N$4639 N$4640 "Straight Waveguide" sch_x=39 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2321 N$4641 N$4642 "Straight Waveguide" sch_x=39 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2322 N$4643 N$4644 "Straight Waveguide" sch_x=39 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2323 N$4645 N$4646 "Straight Waveguide" sch_x=39 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2324 N$4647 N$4648 "Straight Waveguide" sch_x=39 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2325 N$4649 N$4650 "Straight Waveguide" sch_x=37 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2326 N$4651 N$4652 "Straight Waveguide" sch_x=37 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2327 N$4653 N$4654 "Straight Waveguide" sch_x=37 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2328 N$4655 N$4656 "Straight Waveguide" sch_x=37 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2329 N$4657 N$4658 "Straight Waveguide" sch_x=37 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2330 N$4659 N$4660 "Straight Waveguide" sch_x=37 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2331 N$4661 N$4662 "Straight Waveguide" sch_x=35 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2332 N$4663 N$4664 "Straight Waveguide" sch_x=35 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2333 N$4665 N$4666 "Straight Waveguide" sch_x=35 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2334 N$4667 N$4668 "Straight Waveguide" sch_x=35 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2335 N$4669 N$4670 "Straight Waveguide" sch_x=33 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2336 N$4671 N$4672 "Straight Waveguide" sch_x=33 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2337 N$4674 N$4673 "Straight Waveguide" sch_x=45 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2338 N$4676 N$4675 "Straight Waveguide" sch_x=44 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2339 N$4678 N$4677 "Straight Waveguide" sch_x=43 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2340 N$4680 N$4679 "Straight Waveguide" sch_x=42 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2341 N$4682 N$4681 "Straight Waveguide" sch_x=41 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2342 N$4684 N$4683 "Straight Waveguide" sch_x=40 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2343 N$4686 N$4685 "Straight Waveguide" sch_x=39 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2344 N$4688 N$4687 "Straight Waveguide" sch_x=38 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2345 N$4690 N$4689 "Straight Waveguide" sch_x=37 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2346 N$4692 N$4691 "Straight Waveguide" sch_x=36 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2347 N$4694 N$4693 "Straight Waveguide" sch_x=35 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2348 N$4696 N$4695 "Straight Waveguide" sch_x=34 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2349 N$4698 N$4697 "Straight Waveguide" sch_x=33 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2350 N$4700 N$4699 "Straight Waveguide" sch_x=32 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2351 N$4702 N$4701 "Straight Waveguide" sch_x=31 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2352 N$4704 N$4703 "Straight Waveguide" sch_x=31 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2353 N$4706 N$4705 "Straight Waveguide" sch_x=32 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2354 N$4708 N$4707 "Straight Waveguide" sch_x=33 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2355 N$4710 N$4709 "Straight Waveguide" sch_x=34 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2356 N$4712 N$4711 "Straight Waveguide" sch_x=35 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2357 N$4714 N$4713 "Straight Waveguide" sch_x=36 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2358 N$4716 N$4715 "Straight Waveguide" sch_x=37 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2359 N$4718 N$4717 "Straight Waveguide" sch_x=38 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2360 N$4720 N$4719 "Straight Waveguide" sch_x=39 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2361 N$4722 N$4721 "Straight Waveguide" sch_x=40 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2362 N$4724 N$4723 "Straight Waveguide" sch_x=41 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2363 N$4726 N$4725 "Straight Waveguide" sch_x=42 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2364 N$4728 N$4727 "Straight Waveguide" sch_x=43 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2365 N$4730 N$4729 "Straight Waveguide" sch_x=44 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2366 N$4732 N$4731 "Straight Waveguide" sch_x=45 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2367 N$4734 N$4733 "Straight Waveguide" sch_x=46 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2368 N$4736 N$4735 "Straight Waveguide" sch_x=46 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2369 N$4738 N$4737 "Straight Waveguide" sch_x=-125 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2370 N$4740 N$4739 "Straight Waveguide" sch_x=-125 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2371 N$4742 N$4741 "Straight Waveguide" sch_x=-125 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2372 N$4744 N$4743 "Straight Waveguide" sch_x=-125 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2373 N$4746 N$4745 "Straight Waveguide" sch_x=-125 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2374 N$4748 N$4747 "Straight Waveguide" sch_x=-125 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2375 N$4750 N$4749 "Straight Waveguide" sch_x=-125 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2376 N$4752 N$4751 "Straight Waveguide" sch_x=-125 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2377 N$4754 N$4753 "Straight Waveguide" sch_x=-125 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2378 N$4756 N$4755 "Straight Waveguide" sch_x=-125 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2379 N$4758 N$4757 "Straight Waveguide" sch_x=-125 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2380 N$4760 N$4759 "Straight Waveguide" sch_x=-125 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2381 N$4762 N$4761 "Straight Waveguide" sch_x=-125 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2382 N$4764 N$4763 "Straight Waveguide" sch_x=-125 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2383 N$4766 N$4765 "Straight Waveguide" sch_x=-125 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2384 N$4768 N$4767 "Straight Waveguide" sch_x=-125 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2385 N$4770 N$4769 "Straight Waveguide" sch_x=-125 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2386 N$4772 N$4771 "Straight Waveguide" sch_x=-125 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2387 N$4774 N$4773 "Straight Waveguide" sch_x=-125 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2388 N$4776 N$4775 "Straight Waveguide" sch_x=-125 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2389 N$4778 N$4777 "Straight Waveguide" sch_x=-125 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2390 N$4780 N$4779 "Straight Waveguide" sch_x=-125 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2391 N$4782 N$4781 "Straight Waveguide" sch_x=-125 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2392 N$4784 N$4783 "Straight Waveguide" sch_x=-125 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2393 N$4786 N$4785 "Straight Waveguide" sch_x=-125 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2394 N$4788 N$4787 "Straight Waveguide" sch_x=-125 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2395 N$4790 N$4789 "Straight Waveguide" sch_x=-125 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2396 N$4792 N$4791 "Straight Waveguide" sch_x=-125 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2397 N$4794 N$4793 "Straight Waveguide" sch_x=-125 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2398 N$4796 N$4795 "Straight Waveguide" sch_x=-125 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2399 N$4798 N$4797 "Straight Waveguide" sch_x=-125 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2400 N$4800 N$4799 "Straight Waveguide" sch_x=-125 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2401 N$4802 N$4801 "Straight Waveguide" sch_x=-125 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2402 N$4804 N$4803 "Straight Waveguide" sch_x=-125 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2403 N$4806 N$4805 "Straight Waveguide" sch_x=-125 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2404 N$4808 N$4807 "Straight Waveguide" sch_x=-125 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2405 N$4810 N$4809 "Straight Waveguide" sch_x=-125 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2406 N$4812 N$4811 "Straight Waveguide" sch_x=-125 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2407 N$4814 N$4813 "Straight Waveguide" sch_x=-125 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2408 N$4816 N$4815 "Straight Waveguide" sch_x=-125 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2409 N$4818 N$4817 "Straight Waveguide" sch_x=-125 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2410 N$4820 N$4819 "Straight Waveguide" sch_x=-125 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2411 N$4822 N$4821 "Straight Waveguide" sch_x=-125 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2412 N$4824 N$4823 "Straight Waveguide" sch_x=-125 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2413 N$4826 N$4825 "Straight Waveguide" sch_x=-125 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2414 N$4828 N$4827 "Straight Waveguide" sch_x=-125 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2415 N$4830 N$4829 "Straight Waveguide" sch_x=-125 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2416 N$4832 N$4831 "Straight Waveguide" sch_x=-125 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2417 N$4834 N$4833 "Straight Waveguide" sch_x=-125 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2418 N$4836 N$4835 "Straight Waveguide" sch_x=-125 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2419 N$4838 N$4837 "Straight Waveguide" sch_x=-125 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2420 N$4840 N$4839 "Straight Waveguide" sch_x=-125 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2421 N$4842 N$4841 "Straight Waveguide" sch_x=-125 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2422 N$4844 N$4843 "Straight Waveguide" sch_x=-125 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2423 N$4846 N$4845 "Straight Waveguide" sch_x=-125 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2424 N$4848 N$4847 "Straight Waveguide" sch_x=-125 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2425 N$4850 N$4849 "Straight Waveguide" sch_x=-125 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2426 N$4852 N$4851 "Straight Waveguide" sch_x=-125 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2427 N$4854 N$4853 "Straight Waveguide" sch_x=-125 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2428 N$4856 N$4855 "Straight Waveguide" sch_x=-125 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2429 N$4858 N$4857 "Straight Waveguide" sch_x=-125 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2430 N$4860 N$4859 "Straight Waveguide" sch_x=-125 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2431 N$4862 N$4861 "Straight Waveguide" sch_x=-123 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2432 N$4864 N$4863 "Straight Waveguide" sch_x=-123 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2433 N$4866 N$4865 "Straight Waveguide" sch_x=-123 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2434 N$4868 N$4867 "Straight Waveguide" sch_x=-123 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2435 N$4870 N$4869 "Straight Waveguide" sch_x=-123 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2436 N$4872 N$4871 "Straight Waveguide" sch_x=-123 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2437 N$4874 N$4873 "Straight Waveguide" sch_x=-123 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2438 N$4876 N$4875 "Straight Waveguide" sch_x=-123 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2439 N$4878 N$4877 "Straight Waveguide" sch_x=-123 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2440 N$4880 N$4879 "Straight Waveguide" sch_x=-123 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2441 N$4882 N$4881 "Straight Waveguide" sch_x=-123 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2442 N$4884 N$4883 "Straight Waveguide" sch_x=-123 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2443 N$4886 N$4885 "Straight Waveguide" sch_x=-123 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2444 N$4888 N$4887 "Straight Waveguide" sch_x=-123 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2445 N$4890 N$4889 "Straight Waveguide" sch_x=-123 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2446 N$4892 N$4891 "Straight Waveguide" sch_x=-123 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2447 N$4894 N$4893 "Straight Waveguide" sch_x=-123 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2448 N$4896 N$4895 "Straight Waveguide" sch_x=-123 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2449 N$4898 N$4897 "Straight Waveguide" sch_x=-123 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2450 N$4900 N$4899 "Straight Waveguide" sch_x=-123 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2451 N$4902 N$4901 "Straight Waveguide" sch_x=-123 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2452 N$4904 N$4903 "Straight Waveguide" sch_x=-123 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2453 N$4906 N$4905 "Straight Waveguide" sch_x=-123 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2454 N$4908 N$4907 "Straight Waveguide" sch_x=-123 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2455 N$4910 N$4909 "Straight Waveguide" sch_x=-123 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2456 N$4912 N$4911 "Straight Waveguide" sch_x=-123 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2457 N$4914 N$4913 "Straight Waveguide" sch_x=-123 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2458 N$4916 N$4915 "Straight Waveguide" sch_x=-123 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2459 N$4918 N$4917 "Straight Waveguide" sch_x=-123 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2460 N$4920 N$4919 "Straight Waveguide" sch_x=-123 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2461 N$4922 N$4921 "Straight Waveguide" sch_x=-123 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2462 N$4924 N$4923 "Straight Waveguide" sch_x=-123 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2463 N$4926 N$4925 "Straight Waveguide" sch_x=-123 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2464 N$4928 N$4927 "Straight Waveguide" sch_x=-123 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2465 N$4930 N$4929 "Straight Waveguide" sch_x=-123 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2466 N$4932 N$4931 "Straight Waveguide" sch_x=-123 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2467 N$4934 N$4933 "Straight Waveguide" sch_x=-123 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2468 N$4936 N$4935 "Straight Waveguide" sch_x=-123 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2469 N$4938 N$4937 "Straight Waveguide" sch_x=-123 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2470 N$4940 N$4939 "Straight Waveguide" sch_x=-123 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2471 N$4942 N$4941 "Straight Waveguide" sch_x=-123 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2472 N$4944 N$4943 "Straight Waveguide" sch_x=-123 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2473 N$4946 N$4945 "Straight Waveguide" sch_x=-123 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2474 N$4948 N$4947 "Straight Waveguide" sch_x=-123 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2475 N$4950 N$4949 "Straight Waveguide" sch_x=-123 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2476 N$4952 N$4951 "Straight Waveguide" sch_x=-123 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2477 N$4954 N$4953 "Straight Waveguide" sch_x=-123 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2478 N$4956 N$4955 "Straight Waveguide" sch_x=-123 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2479 N$4958 N$4957 "Straight Waveguide" sch_x=-123 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2480 N$4960 N$4959 "Straight Waveguide" sch_x=-123 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2481 N$4962 N$4961 "Straight Waveguide" sch_x=-123 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2482 N$4964 N$4963 "Straight Waveguide" sch_x=-123 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2483 N$4966 N$4965 "Straight Waveguide" sch_x=-123 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2484 N$4968 N$4967 "Straight Waveguide" sch_x=-123 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2485 N$4970 N$4969 "Straight Waveguide" sch_x=-123 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2486 N$4972 N$4971 "Straight Waveguide" sch_x=-123 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2487 N$4974 N$4973 "Straight Waveguide" sch_x=-123 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2488 N$4976 N$4975 "Straight Waveguide" sch_x=-123 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2489 N$4978 N$4977 "Straight Waveguide" sch_x=-123 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2490 N$4980 N$4979 "Straight Waveguide" sch_x=-123 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2491 N$4982 N$4981 "Straight Waveguide" sch_x=-121 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2492 N$4984 N$4983 "Straight Waveguide" sch_x=-121 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2493 N$4986 N$4985 "Straight Waveguide" sch_x=-121 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2494 N$4988 N$4987 "Straight Waveguide" sch_x=-121 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2495 N$4990 N$4989 "Straight Waveguide" sch_x=-121 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2496 N$4992 N$4991 "Straight Waveguide" sch_x=-121 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2497 N$4994 N$4993 "Straight Waveguide" sch_x=-121 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2498 N$4996 N$4995 "Straight Waveguide" sch_x=-121 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2499 N$4998 N$4997 "Straight Waveguide" sch_x=-121 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2500 N$5000 N$4999 "Straight Waveguide" sch_x=-121 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2501 N$5002 N$5001 "Straight Waveguide" sch_x=-121 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2502 N$5004 N$5003 "Straight Waveguide" sch_x=-121 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2503 N$5006 N$5005 "Straight Waveguide" sch_x=-121 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2504 N$5008 N$5007 "Straight Waveguide" sch_x=-121 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2505 N$5010 N$5009 "Straight Waveguide" sch_x=-121 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2506 N$5012 N$5011 "Straight Waveguide" sch_x=-121 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2507 N$5014 N$5013 "Straight Waveguide" sch_x=-121 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2508 N$5016 N$5015 "Straight Waveguide" sch_x=-121 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2509 N$5018 N$5017 "Straight Waveguide" sch_x=-121 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2510 N$5020 N$5019 "Straight Waveguide" sch_x=-121 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2511 N$5022 N$5021 "Straight Waveguide" sch_x=-121 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2512 N$5024 N$5023 "Straight Waveguide" sch_x=-121 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2513 N$5026 N$5025 "Straight Waveguide" sch_x=-121 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2514 N$5028 N$5027 "Straight Waveguide" sch_x=-121 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2515 N$5030 N$5029 "Straight Waveguide" sch_x=-121 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2516 N$5032 N$5031 "Straight Waveguide" sch_x=-121 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2517 N$5034 N$5033 "Straight Waveguide" sch_x=-121 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2518 N$5036 N$5035 "Straight Waveguide" sch_x=-121 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2519 N$5038 N$5037 "Straight Waveguide" sch_x=-121 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2520 N$5040 N$5039 "Straight Waveguide" sch_x=-121 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2521 N$5042 N$5041 "Straight Waveguide" sch_x=-121 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2522 N$5044 N$5043 "Straight Waveguide" sch_x=-121 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2523 N$5046 N$5045 "Straight Waveguide" sch_x=-121 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2524 N$5048 N$5047 "Straight Waveguide" sch_x=-121 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2525 N$5050 N$5049 "Straight Waveguide" sch_x=-121 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2526 N$5052 N$5051 "Straight Waveguide" sch_x=-121 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2527 N$5054 N$5053 "Straight Waveguide" sch_x=-121 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2528 N$5056 N$5055 "Straight Waveguide" sch_x=-121 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2529 N$5058 N$5057 "Straight Waveguide" sch_x=-121 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2530 N$5060 N$5059 "Straight Waveguide" sch_x=-121 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2531 N$5062 N$5061 "Straight Waveguide" sch_x=-121 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2532 N$5064 N$5063 "Straight Waveguide" sch_x=-121 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2533 N$5066 N$5065 "Straight Waveguide" sch_x=-121 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2534 N$5068 N$5067 "Straight Waveguide" sch_x=-121 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2535 N$5070 N$5069 "Straight Waveguide" sch_x=-121 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2536 N$5072 N$5071 "Straight Waveguide" sch_x=-121 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2537 N$5074 N$5073 "Straight Waveguide" sch_x=-121 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2538 N$5076 N$5075 "Straight Waveguide" sch_x=-121 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2539 N$5078 N$5077 "Straight Waveguide" sch_x=-121 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2540 N$5080 N$5079 "Straight Waveguide" sch_x=-121 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2541 N$5082 N$5081 "Straight Waveguide" sch_x=-121 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2542 N$5084 N$5083 "Straight Waveguide" sch_x=-121 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2543 N$5086 N$5085 "Straight Waveguide" sch_x=-121 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2544 N$5088 N$5087 "Straight Waveguide" sch_x=-121 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2545 N$5090 N$5089 "Straight Waveguide" sch_x=-121 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2546 N$5092 N$5091 "Straight Waveguide" sch_x=-121 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2547 N$5094 N$5093 "Straight Waveguide" sch_x=-121 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2548 N$5096 N$5095 "Straight Waveguide" sch_x=-121 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2549 N$5098 N$5097 "Straight Waveguide" sch_x=-119 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2550 N$5100 N$5099 "Straight Waveguide" sch_x=-119 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2551 N$5102 N$5101 "Straight Waveguide" sch_x=-119 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2552 N$5104 N$5103 "Straight Waveguide" sch_x=-119 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2553 N$5106 N$5105 "Straight Waveguide" sch_x=-119 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2554 N$5108 N$5107 "Straight Waveguide" sch_x=-119 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2555 N$5110 N$5109 "Straight Waveguide" sch_x=-119 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2556 N$5112 N$5111 "Straight Waveguide" sch_x=-119 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2557 N$5114 N$5113 "Straight Waveguide" sch_x=-119 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2558 N$5116 N$5115 "Straight Waveguide" sch_x=-119 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2559 N$5118 N$5117 "Straight Waveguide" sch_x=-119 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2560 N$5120 N$5119 "Straight Waveguide" sch_x=-119 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2561 N$5122 N$5121 "Straight Waveguide" sch_x=-119 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2562 N$5124 N$5123 "Straight Waveguide" sch_x=-119 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2563 N$5126 N$5125 "Straight Waveguide" sch_x=-119 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2564 N$5128 N$5127 "Straight Waveguide" sch_x=-119 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2565 N$5130 N$5129 "Straight Waveguide" sch_x=-119 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2566 N$5132 N$5131 "Straight Waveguide" sch_x=-119 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2567 N$5134 N$5133 "Straight Waveguide" sch_x=-119 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2568 N$5136 N$5135 "Straight Waveguide" sch_x=-119 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2569 N$5138 N$5137 "Straight Waveguide" sch_x=-119 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2570 N$5140 N$5139 "Straight Waveguide" sch_x=-119 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2571 N$5142 N$5141 "Straight Waveguide" sch_x=-119 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2572 N$5144 N$5143 "Straight Waveguide" sch_x=-119 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2573 N$5146 N$5145 "Straight Waveguide" sch_x=-119 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2574 N$5148 N$5147 "Straight Waveguide" sch_x=-119 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2575 N$5150 N$5149 "Straight Waveguide" sch_x=-119 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2576 N$5152 N$5151 "Straight Waveguide" sch_x=-119 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2577 N$5154 N$5153 "Straight Waveguide" sch_x=-119 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2578 N$5156 N$5155 "Straight Waveguide" sch_x=-119 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2579 N$5158 N$5157 "Straight Waveguide" sch_x=-119 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2580 N$5160 N$5159 "Straight Waveguide" sch_x=-119 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2581 N$5162 N$5161 "Straight Waveguide" sch_x=-119 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2582 N$5164 N$5163 "Straight Waveguide" sch_x=-119 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2583 N$5166 N$5165 "Straight Waveguide" sch_x=-119 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2584 N$5168 N$5167 "Straight Waveguide" sch_x=-119 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2585 N$5170 N$5169 "Straight Waveguide" sch_x=-119 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2586 N$5172 N$5171 "Straight Waveguide" sch_x=-119 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2587 N$5174 N$5173 "Straight Waveguide" sch_x=-119 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2588 N$5176 N$5175 "Straight Waveguide" sch_x=-119 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2589 N$5178 N$5177 "Straight Waveguide" sch_x=-119 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2590 N$5180 N$5179 "Straight Waveguide" sch_x=-119 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2591 N$5182 N$5181 "Straight Waveguide" sch_x=-119 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2592 N$5184 N$5183 "Straight Waveguide" sch_x=-119 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2593 N$5186 N$5185 "Straight Waveguide" sch_x=-119 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2594 N$5188 N$5187 "Straight Waveguide" sch_x=-119 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2595 N$5190 N$5189 "Straight Waveguide" sch_x=-119 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2596 N$5192 N$5191 "Straight Waveguide" sch_x=-119 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2597 N$5194 N$5193 "Straight Waveguide" sch_x=-119 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2598 N$5196 N$5195 "Straight Waveguide" sch_x=-119 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2599 N$5198 N$5197 "Straight Waveguide" sch_x=-119 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2600 N$5200 N$5199 "Straight Waveguide" sch_x=-119 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2601 N$5202 N$5201 "Straight Waveguide" sch_x=-119 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2602 N$5204 N$5203 "Straight Waveguide" sch_x=-119 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2603 N$5206 N$5205 "Straight Waveguide" sch_x=-119 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2604 N$5208 N$5207 "Straight Waveguide" sch_x=-119 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2605 N$5210 N$5209 "Straight Waveguide" sch_x=-117 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2606 N$5212 N$5211 "Straight Waveguide" sch_x=-117 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2607 N$5214 N$5213 "Straight Waveguide" sch_x=-117 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2608 N$5216 N$5215 "Straight Waveguide" sch_x=-117 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2609 N$5218 N$5217 "Straight Waveguide" sch_x=-117 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2610 N$5220 N$5219 "Straight Waveguide" sch_x=-117 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2611 N$5222 N$5221 "Straight Waveguide" sch_x=-117 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2612 N$5224 N$5223 "Straight Waveguide" sch_x=-117 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2613 N$5226 N$5225 "Straight Waveguide" sch_x=-117 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2614 N$5228 N$5227 "Straight Waveguide" sch_x=-117 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2615 N$5230 N$5229 "Straight Waveguide" sch_x=-117 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2616 N$5232 N$5231 "Straight Waveguide" sch_x=-117 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2617 N$5234 N$5233 "Straight Waveguide" sch_x=-117 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2618 N$5236 N$5235 "Straight Waveguide" sch_x=-117 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2619 N$5238 N$5237 "Straight Waveguide" sch_x=-117 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2620 N$5240 N$5239 "Straight Waveguide" sch_x=-117 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2621 N$5242 N$5241 "Straight Waveguide" sch_x=-117 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2622 N$5244 N$5243 "Straight Waveguide" sch_x=-117 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2623 N$5246 N$5245 "Straight Waveguide" sch_x=-117 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2624 N$5248 N$5247 "Straight Waveguide" sch_x=-117 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2625 N$5250 N$5249 "Straight Waveguide" sch_x=-117 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2626 N$5252 N$5251 "Straight Waveguide" sch_x=-117 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2627 N$5254 N$5253 "Straight Waveguide" sch_x=-117 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2628 N$5256 N$5255 "Straight Waveguide" sch_x=-117 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2629 N$5258 N$5257 "Straight Waveguide" sch_x=-117 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2630 N$5260 N$5259 "Straight Waveguide" sch_x=-117 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2631 N$5262 N$5261 "Straight Waveguide" sch_x=-117 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2632 N$5264 N$5263 "Straight Waveguide" sch_x=-117 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2633 N$5266 N$5265 "Straight Waveguide" sch_x=-117 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2634 N$5268 N$5267 "Straight Waveguide" sch_x=-117 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2635 N$5270 N$5269 "Straight Waveguide" sch_x=-117 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2636 N$5272 N$5271 "Straight Waveguide" sch_x=-117 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2637 N$5274 N$5273 "Straight Waveguide" sch_x=-117 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2638 N$5276 N$5275 "Straight Waveguide" sch_x=-117 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2639 N$5278 N$5277 "Straight Waveguide" sch_x=-117 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2640 N$5280 N$5279 "Straight Waveguide" sch_x=-117 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2641 N$5282 N$5281 "Straight Waveguide" sch_x=-117 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2642 N$5284 N$5283 "Straight Waveguide" sch_x=-117 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2643 N$5286 N$5285 "Straight Waveguide" sch_x=-117 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2644 N$5288 N$5287 "Straight Waveguide" sch_x=-117 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2645 N$5290 N$5289 "Straight Waveguide" sch_x=-117 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2646 N$5292 N$5291 "Straight Waveguide" sch_x=-117 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2647 N$5294 N$5293 "Straight Waveguide" sch_x=-117 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2648 N$5296 N$5295 "Straight Waveguide" sch_x=-117 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2649 N$5298 N$5297 "Straight Waveguide" sch_x=-117 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2650 N$5300 N$5299 "Straight Waveguide" sch_x=-117 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2651 N$5302 N$5301 "Straight Waveguide" sch_x=-117 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2652 N$5304 N$5303 "Straight Waveguide" sch_x=-117 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2653 N$5306 N$5305 "Straight Waveguide" sch_x=-117 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2654 N$5308 N$5307 "Straight Waveguide" sch_x=-117 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2655 N$5310 N$5309 "Straight Waveguide" sch_x=-117 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2656 N$5312 N$5311 "Straight Waveguide" sch_x=-117 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2657 N$5314 N$5313 "Straight Waveguide" sch_x=-117 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2658 N$5316 N$5315 "Straight Waveguide" sch_x=-117 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2659 N$5318 N$5317 "Straight Waveguide" sch_x=-115 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2660 N$5320 N$5319 "Straight Waveguide" sch_x=-115 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2661 N$5322 N$5321 "Straight Waveguide" sch_x=-115 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2662 N$5324 N$5323 "Straight Waveguide" sch_x=-115 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2663 N$5326 N$5325 "Straight Waveguide" sch_x=-115 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2664 N$5328 N$5327 "Straight Waveguide" sch_x=-115 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2665 N$5330 N$5329 "Straight Waveguide" sch_x=-115 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2666 N$5332 N$5331 "Straight Waveguide" sch_x=-115 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2667 N$5334 N$5333 "Straight Waveguide" sch_x=-115 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2668 N$5336 N$5335 "Straight Waveguide" sch_x=-115 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2669 N$5338 N$5337 "Straight Waveguide" sch_x=-115 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2670 N$5340 N$5339 "Straight Waveguide" sch_x=-115 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2671 N$5342 N$5341 "Straight Waveguide" sch_x=-115 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2672 N$5344 N$5343 "Straight Waveguide" sch_x=-115 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2673 N$5346 N$5345 "Straight Waveguide" sch_x=-115 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2674 N$5348 N$5347 "Straight Waveguide" sch_x=-115 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2675 N$5350 N$5349 "Straight Waveguide" sch_x=-115 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2676 N$5352 N$5351 "Straight Waveguide" sch_x=-115 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2677 N$5354 N$5353 "Straight Waveguide" sch_x=-115 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2678 N$5356 N$5355 "Straight Waveguide" sch_x=-115 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2679 N$5358 N$5357 "Straight Waveguide" sch_x=-115 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2680 N$5360 N$5359 "Straight Waveguide" sch_x=-115 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2681 N$5362 N$5361 "Straight Waveguide" sch_x=-115 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2682 N$5364 N$5363 "Straight Waveguide" sch_x=-115 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2683 N$5366 N$5365 "Straight Waveguide" sch_x=-115 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2684 N$5368 N$5367 "Straight Waveguide" sch_x=-115 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2685 N$5370 N$5369 "Straight Waveguide" sch_x=-115 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2686 N$5372 N$5371 "Straight Waveguide" sch_x=-115 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2687 N$5374 N$5373 "Straight Waveguide" sch_x=-115 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2688 N$5376 N$5375 "Straight Waveguide" sch_x=-115 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2689 N$5378 N$5377 "Straight Waveguide" sch_x=-115 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2690 N$5380 N$5379 "Straight Waveguide" sch_x=-115 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2691 N$5382 N$5381 "Straight Waveguide" sch_x=-115 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2692 N$5384 N$5383 "Straight Waveguide" sch_x=-115 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2693 N$5386 N$5385 "Straight Waveguide" sch_x=-115 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2694 N$5388 N$5387 "Straight Waveguide" sch_x=-115 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2695 N$5390 N$5389 "Straight Waveguide" sch_x=-115 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2696 N$5392 N$5391 "Straight Waveguide" sch_x=-115 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2697 N$5394 N$5393 "Straight Waveguide" sch_x=-115 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2698 N$5396 N$5395 "Straight Waveguide" sch_x=-115 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2699 N$5398 N$5397 "Straight Waveguide" sch_x=-115 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2700 N$5400 N$5399 "Straight Waveguide" sch_x=-115 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2701 N$5402 N$5401 "Straight Waveguide" sch_x=-115 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2702 N$5404 N$5403 "Straight Waveguide" sch_x=-115 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2703 N$5406 N$5405 "Straight Waveguide" sch_x=-115 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2704 N$5408 N$5407 "Straight Waveguide" sch_x=-115 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2705 N$5410 N$5409 "Straight Waveguide" sch_x=-115 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2706 N$5412 N$5411 "Straight Waveguide" sch_x=-115 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2707 N$5414 N$5413 "Straight Waveguide" sch_x=-115 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2708 N$5416 N$5415 "Straight Waveguide" sch_x=-115 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2709 N$5418 N$5417 "Straight Waveguide" sch_x=-115 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2710 N$5420 N$5419 "Straight Waveguide" sch_x=-115 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2711 N$5422 N$5421 "Straight Waveguide" sch_x=-113 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2712 N$5424 N$5423 "Straight Waveguide" sch_x=-113 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2713 N$5426 N$5425 "Straight Waveguide" sch_x=-113 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2714 N$5428 N$5427 "Straight Waveguide" sch_x=-113 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2715 N$5430 N$5429 "Straight Waveguide" sch_x=-113 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2716 N$5432 N$5431 "Straight Waveguide" sch_x=-113 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2717 N$5434 N$5433 "Straight Waveguide" sch_x=-113 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2718 N$5436 N$5435 "Straight Waveguide" sch_x=-113 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2719 N$5438 N$5437 "Straight Waveguide" sch_x=-113 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2720 N$5440 N$5439 "Straight Waveguide" sch_x=-113 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2721 N$5442 N$5441 "Straight Waveguide" sch_x=-113 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2722 N$5444 N$5443 "Straight Waveguide" sch_x=-113 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2723 N$5446 N$5445 "Straight Waveguide" sch_x=-113 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2724 N$5448 N$5447 "Straight Waveguide" sch_x=-113 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2725 N$5450 N$5449 "Straight Waveguide" sch_x=-113 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2726 N$5452 N$5451 "Straight Waveguide" sch_x=-113 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2727 N$5454 N$5453 "Straight Waveguide" sch_x=-113 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2728 N$5456 N$5455 "Straight Waveguide" sch_x=-113 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2729 N$5458 N$5457 "Straight Waveguide" sch_x=-113 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2730 N$5460 N$5459 "Straight Waveguide" sch_x=-113 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2731 N$5462 N$5461 "Straight Waveguide" sch_x=-113 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2732 N$5464 N$5463 "Straight Waveguide" sch_x=-113 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2733 N$5466 N$5465 "Straight Waveguide" sch_x=-113 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2734 N$5468 N$5467 "Straight Waveguide" sch_x=-113 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2735 N$5470 N$5469 "Straight Waveguide" sch_x=-113 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2736 N$5472 N$5471 "Straight Waveguide" sch_x=-113 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2737 N$5474 N$5473 "Straight Waveguide" sch_x=-113 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2738 N$5476 N$5475 "Straight Waveguide" sch_x=-113 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2739 N$5478 N$5477 "Straight Waveguide" sch_x=-113 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2740 N$5480 N$5479 "Straight Waveguide" sch_x=-113 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2741 N$5482 N$5481 "Straight Waveguide" sch_x=-113 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2742 N$5484 N$5483 "Straight Waveguide" sch_x=-113 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2743 N$5486 N$5485 "Straight Waveguide" sch_x=-113 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2744 N$5488 N$5487 "Straight Waveguide" sch_x=-113 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2745 N$5490 N$5489 "Straight Waveguide" sch_x=-113 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2746 N$5492 N$5491 "Straight Waveguide" sch_x=-113 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2747 N$5494 N$5493 "Straight Waveguide" sch_x=-113 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2748 N$5496 N$5495 "Straight Waveguide" sch_x=-113 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2749 N$5498 N$5497 "Straight Waveguide" sch_x=-113 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2750 N$5500 N$5499 "Straight Waveguide" sch_x=-113 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2751 N$5502 N$5501 "Straight Waveguide" sch_x=-113 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2752 N$5504 N$5503 "Straight Waveguide" sch_x=-113 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2753 N$5506 N$5505 "Straight Waveguide" sch_x=-113 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2754 N$5508 N$5507 "Straight Waveguide" sch_x=-113 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2755 N$5510 N$5509 "Straight Waveguide" sch_x=-113 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2756 N$5512 N$5511 "Straight Waveguide" sch_x=-113 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2757 N$5514 N$5513 "Straight Waveguide" sch_x=-113 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2758 N$5516 N$5515 "Straight Waveguide" sch_x=-113 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2759 N$5518 N$5517 "Straight Waveguide" sch_x=-113 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2760 N$5520 N$5519 "Straight Waveguide" sch_x=-113 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2761 N$5522 N$5521 "Straight Waveguide" sch_x=-111 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2762 N$5524 N$5523 "Straight Waveguide" sch_x=-111 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2763 N$5526 N$5525 "Straight Waveguide" sch_x=-111 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2764 N$5528 N$5527 "Straight Waveguide" sch_x=-111 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2765 N$5530 N$5529 "Straight Waveguide" sch_x=-111 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2766 N$5532 N$5531 "Straight Waveguide" sch_x=-111 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2767 N$5534 N$5533 "Straight Waveguide" sch_x=-111 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2768 N$5536 N$5535 "Straight Waveguide" sch_x=-111 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2769 N$5538 N$5537 "Straight Waveguide" sch_x=-111 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2770 N$5540 N$5539 "Straight Waveguide" sch_x=-111 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2771 N$5542 N$5541 "Straight Waveguide" sch_x=-111 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2772 N$5544 N$5543 "Straight Waveguide" sch_x=-111 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2773 N$5546 N$5545 "Straight Waveguide" sch_x=-111 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2774 N$5548 N$5547 "Straight Waveguide" sch_x=-111 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2775 N$5550 N$5549 "Straight Waveguide" sch_x=-111 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2776 N$5552 N$5551 "Straight Waveguide" sch_x=-111 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2777 N$5554 N$5553 "Straight Waveguide" sch_x=-111 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2778 N$5556 N$5555 "Straight Waveguide" sch_x=-111 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2779 N$5558 N$5557 "Straight Waveguide" sch_x=-111 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2780 N$5560 N$5559 "Straight Waveguide" sch_x=-111 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2781 N$5562 N$5561 "Straight Waveguide" sch_x=-111 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2782 N$5564 N$5563 "Straight Waveguide" sch_x=-111 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2783 N$5566 N$5565 "Straight Waveguide" sch_x=-111 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2784 N$5568 N$5567 "Straight Waveguide" sch_x=-111 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2785 N$5570 N$5569 "Straight Waveguide" sch_x=-111 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2786 N$5572 N$5571 "Straight Waveguide" sch_x=-111 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2787 N$5574 N$5573 "Straight Waveguide" sch_x=-111 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2788 N$5576 N$5575 "Straight Waveguide" sch_x=-111 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2789 N$5578 N$5577 "Straight Waveguide" sch_x=-111 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2790 N$5580 N$5579 "Straight Waveguide" sch_x=-111 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2791 N$5582 N$5581 "Straight Waveguide" sch_x=-111 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2792 N$5584 N$5583 "Straight Waveguide" sch_x=-111 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2793 N$5586 N$5585 "Straight Waveguide" sch_x=-111 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2794 N$5588 N$5587 "Straight Waveguide" sch_x=-111 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2795 N$5590 N$5589 "Straight Waveguide" sch_x=-111 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2796 N$5592 N$5591 "Straight Waveguide" sch_x=-111 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2797 N$5594 N$5593 "Straight Waveguide" sch_x=-111 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2798 N$5596 N$5595 "Straight Waveguide" sch_x=-111 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2799 N$5598 N$5597 "Straight Waveguide" sch_x=-111 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2800 N$5600 N$5599 "Straight Waveguide" sch_x=-111 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2801 N$5602 N$5601 "Straight Waveguide" sch_x=-111 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2802 N$5604 N$5603 "Straight Waveguide" sch_x=-111 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2803 N$5606 N$5605 "Straight Waveguide" sch_x=-111 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2804 N$5608 N$5607 "Straight Waveguide" sch_x=-111 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2805 N$5610 N$5609 "Straight Waveguide" sch_x=-111 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2806 N$5612 N$5611 "Straight Waveguide" sch_x=-111 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2807 N$5614 N$5613 "Straight Waveguide" sch_x=-111 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2808 N$5616 N$5615 "Straight Waveguide" sch_x=-111 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2809 N$5618 N$5617 "Straight Waveguide" sch_x=-109 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2810 N$5620 N$5619 "Straight Waveguide" sch_x=-109 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2811 N$5622 N$5621 "Straight Waveguide" sch_x=-109 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2812 N$5624 N$5623 "Straight Waveguide" sch_x=-109 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2813 N$5626 N$5625 "Straight Waveguide" sch_x=-109 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2814 N$5628 N$5627 "Straight Waveguide" sch_x=-109 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2815 N$5630 N$5629 "Straight Waveguide" sch_x=-109 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2816 N$5632 N$5631 "Straight Waveguide" sch_x=-109 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2817 N$5634 N$5633 "Straight Waveguide" sch_x=-109 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2818 N$5636 N$5635 "Straight Waveguide" sch_x=-109 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2819 N$5638 N$5637 "Straight Waveguide" sch_x=-109 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2820 N$5640 N$5639 "Straight Waveguide" sch_x=-109 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2821 N$5642 N$5641 "Straight Waveguide" sch_x=-109 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2822 N$5644 N$5643 "Straight Waveguide" sch_x=-109 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2823 N$5646 N$5645 "Straight Waveguide" sch_x=-109 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2824 N$5648 N$5647 "Straight Waveguide" sch_x=-109 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2825 N$5650 N$5649 "Straight Waveguide" sch_x=-109 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2826 N$5652 N$5651 "Straight Waveguide" sch_x=-109 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2827 N$5654 N$5653 "Straight Waveguide" sch_x=-109 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2828 N$5656 N$5655 "Straight Waveguide" sch_x=-109 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2829 N$5658 N$5657 "Straight Waveguide" sch_x=-109 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2830 N$5660 N$5659 "Straight Waveguide" sch_x=-109 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2831 N$5662 N$5661 "Straight Waveguide" sch_x=-109 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2832 N$5664 N$5663 "Straight Waveguide" sch_x=-109 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2833 N$5666 N$5665 "Straight Waveguide" sch_x=-109 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2834 N$5668 N$5667 "Straight Waveguide" sch_x=-109 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2835 N$5670 N$5669 "Straight Waveguide" sch_x=-109 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2836 N$5672 N$5671 "Straight Waveguide" sch_x=-109 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2837 N$5674 N$5673 "Straight Waveguide" sch_x=-109 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2838 N$5676 N$5675 "Straight Waveguide" sch_x=-109 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2839 N$5678 N$5677 "Straight Waveguide" sch_x=-109 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2840 N$5680 N$5679 "Straight Waveguide" sch_x=-109 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2841 N$5682 N$5681 "Straight Waveguide" sch_x=-109 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2842 N$5684 N$5683 "Straight Waveguide" sch_x=-109 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2843 N$5686 N$5685 "Straight Waveguide" sch_x=-109 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2844 N$5688 N$5687 "Straight Waveguide" sch_x=-109 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2845 N$5690 N$5689 "Straight Waveguide" sch_x=-109 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2846 N$5692 N$5691 "Straight Waveguide" sch_x=-109 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2847 N$5694 N$5693 "Straight Waveguide" sch_x=-109 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2848 N$5696 N$5695 "Straight Waveguide" sch_x=-109 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2849 N$5698 N$5697 "Straight Waveguide" sch_x=-109 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2850 N$5700 N$5699 "Straight Waveguide" sch_x=-109 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2851 N$5702 N$5701 "Straight Waveguide" sch_x=-109 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2852 N$5704 N$5703 "Straight Waveguide" sch_x=-109 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2853 N$5706 N$5705 "Straight Waveguide" sch_x=-109 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2854 N$5708 N$5707 "Straight Waveguide" sch_x=-109 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2855 N$5710 N$5709 "Straight Waveguide" sch_x=-107 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2856 N$5712 N$5711 "Straight Waveguide" sch_x=-107 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2857 N$5714 N$5713 "Straight Waveguide" sch_x=-107 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2858 N$5716 N$5715 "Straight Waveguide" sch_x=-107 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2859 N$5718 N$5717 "Straight Waveguide" sch_x=-107 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2860 N$5720 N$5719 "Straight Waveguide" sch_x=-107 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2861 N$5722 N$5721 "Straight Waveguide" sch_x=-107 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2862 N$5724 N$5723 "Straight Waveguide" sch_x=-107 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2863 N$5726 N$5725 "Straight Waveguide" sch_x=-107 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2864 N$5728 N$5727 "Straight Waveguide" sch_x=-107 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2865 N$5730 N$5729 "Straight Waveguide" sch_x=-107 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2866 N$5732 N$5731 "Straight Waveguide" sch_x=-107 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2867 N$5734 N$5733 "Straight Waveguide" sch_x=-107 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2868 N$5736 N$5735 "Straight Waveguide" sch_x=-107 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2869 N$5738 N$5737 "Straight Waveguide" sch_x=-107 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2870 N$5740 N$5739 "Straight Waveguide" sch_x=-107 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2871 N$5742 N$5741 "Straight Waveguide" sch_x=-107 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2872 N$5744 N$5743 "Straight Waveguide" sch_x=-107 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2873 N$5746 N$5745 "Straight Waveguide" sch_x=-107 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2874 N$5748 N$5747 "Straight Waveguide" sch_x=-107 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2875 N$5750 N$5749 "Straight Waveguide" sch_x=-107 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2876 N$5752 N$5751 "Straight Waveguide" sch_x=-107 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2877 N$5754 N$5753 "Straight Waveguide" sch_x=-107 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2878 N$5756 N$5755 "Straight Waveguide" sch_x=-107 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2879 N$5758 N$5757 "Straight Waveguide" sch_x=-107 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2880 N$5760 N$5759 "Straight Waveguide" sch_x=-107 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2881 N$5762 N$5761 "Straight Waveguide" sch_x=-107 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2882 N$5764 N$5763 "Straight Waveguide" sch_x=-107 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2883 N$5766 N$5765 "Straight Waveguide" sch_x=-107 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2884 N$5768 N$5767 "Straight Waveguide" sch_x=-107 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2885 N$5770 N$5769 "Straight Waveguide" sch_x=-107 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2886 N$5772 N$5771 "Straight Waveguide" sch_x=-107 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2887 N$5774 N$5773 "Straight Waveguide" sch_x=-107 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2888 N$5776 N$5775 "Straight Waveguide" sch_x=-107 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2889 N$5778 N$5777 "Straight Waveguide" sch_x=-107 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2890 N$5780 N$5779 "Straight Waveguide" sch_x=-107 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2891 N$5782 N$5781 "Straight Waveguide" sch_x=-107 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2892 N$5784 N$5783 "Straight Waveguide" sch_x=-107 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2893 N$5786 N$5785 "Straight Waveguide" sch_x=-107 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2894 N$5788 N$5787 "Straight Waveguide" sch_x=-107 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2895 N$5790 N$5789 "Straight Waveguide" sch_x=-107 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2896 N$5792 N$5791 "Straight Waveguide" sch_x=-107 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2897 N$5794 N$5793 "Straight Waveguide" sch_x=-107 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2898 N$5796 N$5795 "Straight Waveguide" sch_x=-107 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2899 N$5798 N$5797 "Straight Waveguide" sch_x=-105 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2900 N$5800 N$5799 "Straight Waveguide" sch_x=-105 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2901 N$5802 N$5801 "Straight Waveguide" sch_x=-105 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2902 N$5804 N$5803 "Straight Waveguide" sch_x=-105 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2903 N$5806 N$5805 "Straight Waveguide" sch_x=-105 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2904 N$5808 N$5807 "Straight Waveguide" sch_x=-105 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2905 N$5810 N$5809 "Straight Waveguide" sch_x=-105 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2906 N$5812 N$5811 "Straight Waveguide" sch_x=-105 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2907 N$5814 N$5813 "Straight Waveguide" sch_x=-105 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2908 N$5816 N$5815 "Straight Waveguide" sch_x=-105 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2909 N$5818 N$5817 "Straight Waveguide" sch_x=-105 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2910 N$5820 N$5819 "Straight Waveguide" sch_x=-105 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2911 N$5822 N$5821 "Straight Waveguide" sch_x=-105 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2912 N$5824 N$5823 "Straight Waveguide" sch_x=-105 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2913 N$5826 N$5825 "Straight Waveguide" sch_x=-105 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2914 N$5828 N$5827 "Straight Waveguide" sch_x=-105 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2915 N$5830 N$5829 "Straight Waveguide" sch_x=-105 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2916 N$5832 N$5831 "Straight Waveguide" sch_x=-105 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2917 N$5834 N$5833 "Straight Waveguide" sch_x=-105 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2918 N$5836 N$5835 "Straight Waveguide" sch_x=-105 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2919 N$5838 N$5837 "Straight Waveguide" sch_x=-105 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2920 N$5840 N$5839 "Straight Waveguide" sch_x=-105 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2921 N$5842 N$5841 "Straight Waveguide" sch_x=-105 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2922 N$5844 N$5843 "Straight Waveguide" sch_x=-105 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2923 N$5846 N$5845 "Straight Waveguide" sch_x=-105 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2924 N$5848 N$5847 "Straight Waveguide" sch_x=-105 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2925 N$5850 N$5849 "Straight Waveguide" sch_x=-105 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2926 N$5852 N$5851 "Straight Waveguide" sch_x=-105 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2927 N$5854 N$5853 "Straight Waveguide" sch_x=-105 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2928 N$5856 N$5855 "Straight Waveguide" sch_x=-105 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2929 N$5858 N$5857 "Straight Waveguide" sch_x=-105 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2930 N$5860 N$5859 "Straight Waveguide" sch_x=-105 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2931 N$5862 N$5861 "Straight Waveguide" sch_x=-105 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2932 N$5864 N$5863 "Straight Waveguide" sch_x=-105 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2933 N$5866 N$5865 "Straight Waveguide" sch_x=-105 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2934 N$5868 N$5867 "Straight Waveguide" sch_x=-105 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2935 N$5870 N$5869 "Straight Waveguide" sch_x=-105 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2936 N$5872 N$5871 "Straight Waveguide" sch_x=-105 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2937 N$5874 N$5873 "Straight Waveguide" sch_x=-105 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2938 N$5876 N$5875 "Straight Waveguide" sch_x=-105 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2939 N$5878 N$5877 "Straight Waveguide" sch_x=-105 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2940 N$5880 N$5879 "Straight Waveguide" sch_x=-105 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2941 N$5882 N$5881 "Straight Waveguide" sch_x=-103 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2942 N$5884 N$5883 "Straight Waveguide" sch_x=-103 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2943 N$5886 N$5885 "Straight Waveguide" sch_x=-103 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2944 N$5888 N$5887 "Straight Waveguide" sch_x=-103 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2945 N$5890 N$5889 "Straight Waveguide" sch_x=-103 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2946 N$5892 N$5891 "Straight Waveguide" sch_x=-103 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2947 N$5894 N$5893 "Straight Waveguide" sch_x=-103 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2948 N$5896 N$5895 "Straight Waveguide" sch_x=-103 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2949 N$5898 N$5897 "Straight Waveguide" sch_x=-103 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2950 N$5900 N$5899 "Straight Waveguide" sch_x=-103 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2951 N$5902 N$5901 "Straight Waveguide" sch_x=-103 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2952 N$5904 N$5903 "Straight Waveguide" sch_x=-103 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2953 N$5906 N$5905 "Straight Waveguide" sch_x=-103 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2954 N$5908 N$5907 "Straight Waveguide" sch_x=-103 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2955 N$5910 N$5909 "Straight Waveguide" sch_x=-103 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2956 N$5912 N$5911 "Straight Waveguide" sch_x=-103 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2957 N$5914 N$5913 "Straight Waveguide" sch_x=-103 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2958 N$5916 N$5915 "Straight Waveguide" sch_x=-103 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2959 N$5918 N$5917 "Straight Waveguide" sch_x=-103 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2960 N$5920 N$5919 "Straight Waveguide" sch_x=-103 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2961 N$5922 N$5921 "Straight Waveguide" sch_x=-103 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2962 N$5924 N$5923 "Straight Waveguide" sch_x=-103 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2963 N$5926 N$5925 "Straight Waveguide" sch_x=-103 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2964 N$5928 N$5927 "Straight Waveguide" sch_x=-103 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2965 N$5930 N$5929 "Straight Waveguide" sch_x=-103 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2966 N$5932 N$5931 "Straight Waveguide" sch_x=-103 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2967 N$5934 N$5933 "Straight Waveguide" sch_x=-103 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2968 N$5936 N$5935 "Straight Waveguide" sch_x=-103 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2969 N$5938 N$5937 "Straight Waveguide" sch_x=-103 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2970 N$5940 N$5939 "Straight Waveguide" sch_x=-103 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2971 N$5942 N$5941 "Straight Waveguide" sch_x=-103 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2972 N$5944 N$5943 "Straight Waveguide" sch_x=-103 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2973 N$5946 N$5945 "Straight Waveguide" sch_x=-103 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2974 N$5948 N$5947 "Straight Waveguide" sch_x=-103 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2975 N$5950 N$5949 "Straight Waveguide" sch_x=-103 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2976 N$5952 N$5951 "Straight Waveguide" sch_x=-103 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2977 N$5954 N$5953 "Straight Waveguide" sch_x=-103 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2978 N$5956 N$5955 "Straight Waveguide" sch_x=-103 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2979 N$5958 N$5957 "Straight Waveguide" sch_x=-103 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2980 N$5960 N$5959 "Straight Waveguide" sch_x=-103 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2981 N$5962 N$5961 "Straight Waveguide" sch_x=-101 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2982 N$5964 N$5963 "Straight Waveguide" sch_x=-101 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2983 N$5966 N$5965 "Straight Waveguide" sch_x=-101 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2984 N$5968 N$5967 "Straight Waveguide" sch_x=-101 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2985 N$5970 N$5969 "Straight Waveguide" sch_x=-101 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2986 N$5972 N$5971 "Straight Waveguide" sch_x=-101 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2987 N$5974 N$5973 "Straight Waveguide" sch_x=-101 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2988 N$5976 N$5975 "Straight Waveguide" sch_x=-101 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2989 N$5978 N$5977 "Straight Waveguide" sch_x=-101 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2990 N$5980 N$5979 "Straight Waveguide" sch_x=-101 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2991 N$5982 N$5981 "Straight Waveguide" sch_x=-101 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2992 N$5984 N$5983 "Straight Waveguide" sch_x=-101 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2993 N$5986 N$5985 "Straight Waveguide" sch_x=-101 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2994 N$5988 N$5987 "Straight Waveguide" sch_x=-101 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2995 N$5990 N$5989 "Straight Waveguide" sch_x=-101 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2996 N$5992 N$5991 "Straight Waveguide" sch_x=-101 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2997 N$5994 N$5993 "Straight Waveguide" sch_x=-101 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2998 N$5996 N$5995 "Straight Waveguide" sch_x=-101 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W2999 N$5998 N$5997 "Straight Waveguide" sch_x=-101 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3000 N$6000 N$5999 "Straight Waveguide" sch_x=-101 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3001 N$6002 N$6001 "Straight Waveguide" sch_x=-101 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3002 N$6004 N$6003 "Straight Waveguide" sch_x=-101 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3003 N$6006 N$6005 "Straight Waveguide" sch_x=-101 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3004 N$6008 N$6007 "Straight Waveguide" sch_x=-101 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3005 N$6010 N$6009 "Straight Waveguide" sch_x=-101 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3006 N$6012 N$6011 "Straight Waveguide" sch_x=-101 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3007 N$6014 N$6013 "Straight Waveguide" sch_x=-101 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3008 N$6016 N$6015 "Straight Waveguide" sch_x=-101 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3009 N$6018 N$6017 "Straight Waveguide" sch_x=-101 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3010 N$6020 N$6019 "Straight Waveguide" sch_x=-101 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3011 N$6022 N$6021 "Straight Waveguide" sch_x=-101 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3012 N$6024 N$6023 "Straight Waveguide" sch_x=-101 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3013 N$6026 N$6025 "Straight Waveguide" sch_x=-101 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3014 N$6028 N$6027 "Straight Waveguide" sch_x=-101 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3015 N$6030 N$6029 "Straight Waveguide" sch_x=-101 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3016 N$6032 N$6031 "Straight Waveguide" sch_x=-101 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3017 N$6034 N$6033 "Straight Waveguide" sch_x=-101 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3018 N$6036 N$6035 "Straight Waveguide" sch_x=-101 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3019 N$6038 N$6037 "Straight Waveguide" sch_x=-99 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3020 N$6040 N$6039 "Straight Waveguide" sch_x=-99 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3021 N$6042 N$6041 "Straight Waveguide" sch_x=-99 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3022 N$6044 N$6043 "Straight Waveguide" sch_x=-99 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3023 N$6046 N$6045 "Straight Waveguide" sch_x=-99 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3024 N$6048 N$6047 "Straight Waveguide" sch_x=-99 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3025 N$6050 N$6049 "Straight Waveguide" sch_x=-99 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3026 N$6052 N$6051 "Straight Waveguide" sch_x=-99 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3027 N$6054 N$6053 "Straight Waveguide" sch_x=-99 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3028 N$6056 N$6055 "Straight Waveguide" sch_x=-99 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3029 N$6058 N$6057 "Straight Waveguide" sch_x=-99 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3030 N$6060 N$6059 "Straight Waveguide" sch_x=-99 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3031 N$6062 N$6061 "Straight Waveguide" sch_x=-99 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3032 N$6064 N$6063 "Straight Waveguide" sch_x=-99 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3033 N$6066 N$6065 "Straight Waveguide" sch_x=-99 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3034 N$6068 N$6067 "Straight Waveguide" sch_x=-99 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3035 N$6070 N$6069 "Straight Waveguide" sch_x=-99 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3036 N$6072 N$6071 "Straight Waveguide" sch_x=-99 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3037 N$6074 N$6073 "Straight Waveguide" sch_x=-99 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3038 N$6076 N$6075 "Straight Waveguide" sch_x=-99 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3039 N$6078 N$6077 "Straight Waveguide" sch_x=-99 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3040 N$6080 N$6079 "Straight Waveguide" sch_x=-99 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3041 N$6082 N$6081 "Straight Waveguide" sch_x=-99 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3042 N$6084 N$6083 "Straight Waveguide" sch_x=-99 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3043 N$6086 N$6085 "Straight Waveguide" sch_x=-99 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3044 N$6088 N$6087 "Straight Waveguide" sch_x=-99 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3045 N$6090 N$6089 "Straight Waveguide" sch_x=-99 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3046 N$6092 N$6091 "Straight Waveguide" sch_x=-99 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3047 N$6094 N$6093 "Straight Waveguide" sch_x=-99 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3048 N$6096 N$6095 "Straight Waveguide" sch_x=-99 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3049 N$6098 N$6097 "Straight Waveguide" sch_x=-99 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3050 N$6100 N$6099 "Straight Waveguide" sch_x=-99 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3051 N$6102 N$6101 "Straight Waveguide" sch_x=-99 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3052 N$6104 N$6103 "Straight Waveguide" sch_x=-99 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3053 N$6106 N$6105 "Straight Waveguide" sch_x=-99 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3054 N$6108 N$6107 "Straight Waveguide" sch_x=-99 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3055 N$6110 N$6109 "Straight Waveguide" sch_x=-97 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3056 N$6112 N$6111 "Straight Waveguide" sch_x=-97 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3057 N$6114 N$6113 "Straight Waveguide" sch_x=-97 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3058 N$6116 N$6115 "Straight Waveguide" sch_x=-97 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3059 N$6118 N$6117 "Straight Waveguide" sch_x=-97 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3060 N$6120 N$6119 "Straight Waveguide" sch_x=-97 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3061 N$6122 N$6121 "Straight Waveguide" sch_x=-97 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3062 N$6124 N$6123 "Straight Waveguide" sch_x=-97 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3063 N$6126 N$6125 "Straight Waveguide" sch_x=-97 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3064 N$6128 N$6127 "Straight Waveguide" sch_x=-97 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3065 N$6130 N$6129 "Straight Waveguide" sch_x=-97 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3066 N$6132 N$6131 "Straight Waveguide" sch_x=-97 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3067 N$6134 N$6133 "Straight Waveguide" sch_x=-97 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3068 N$6136 N$6135 "Straight Waveguide" sch_x=-97 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3069 N$6138 N$6137 "Straight Waveguide" sch_x=-97 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3070 N$6140 N$6139 "Straight Waveguide" sch_x=-97 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3071 N$6142 N$6141 "Straight Waveguide" sch_x=-97 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3072 N$6144 N$6143 "Straight Waveguide" sch_x=-97 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3073 N$6146 N$6145 "Straight Waveguide" sch_x=-97 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3074 N$6148 N$6147 "Straight Waveguide" sch_x=-97 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3075 N$6150 N$6149 "Straight Waveguide" sch_x=-97 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3076 N$6152 N$6151 "Straight Waveguide" sch_x=-97 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3077 N$6154 N$6153 "Straight Waveguide" sch_x=-97 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3078 N$6156 N$6155 "Straight Waveguide" sch_x=-97 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3079 N$6158 N$6157 "Straight Waveguide" sch_x=-97 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3080 N$6160 N$6159 "Straight Waveguide" sch_x=-97 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3081 N$6162 N$6161 "Straight Waveguide" sch_x=-97 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3082 N$6164 N$6163 "Straight Waveguide" sch_x=-97 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3083 N$6166 N$6165 "Straight Waveguide" sch_x=-97 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3084 N$6168 N$6167 "Straight Waveguide" sch_x=-97 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3085 N$6170 N$6169 "Straight Waveguide" sch_x=-97 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3086 N$6172 N$6171 "Straight Waveguide" sch_x=-97 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3087 N$6174 N$6173 "Straight Waveguide" sch_x=-97 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3088 N$6176 N$6175 "Straight Waveguide" sch_x=-97 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3089 N$6178 N$6177 "Straight Waveguide" sch_x=-95 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3090 N$6180 N$6179 "Straight Waveguide" sch_x=-95 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3091 N$6182 N$6181 "Straight Waveguide" sch_x=-95 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3092 N$6184 N$6183 "Straight Waveguide" sch_x=-95 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3093 N$6186 N$6185 "Straight Waveguide" sch_x=-95 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3094 N$6188 N$6187 "Straight Waveguide" sch_x=-95 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3095 N$6190 N$6189 "Straight Waveguide" sch_x=-95 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3096 N$6192 N$6191 "Straight Waveguide" sch_x=-95 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3097 N$6194 N$6193 "Straight Waveguide" sch_x=-95 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3098 N$6196 N$6195 "Straight Waveguide" sch_x=-95 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3099 N$6198 N$6197 "Straight Waveguide" sch_x=-95 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3100 N$6200 N$6199 "Straight Waveguide" sch_x=-95 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3101 N$6202 N$6201 "Straight Waveguide" sch_x=-95 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3102 N$6204 N$6203 "Straight Waveguide" sch_x=-95 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3103 N$6206 N$6205 "Straight Waveguide" sch_x=-95 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3104 N$6208 N$6207 "Straight Waveguide" sch_x=-95 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3105 N$6210 N$6209 "Straight Waveguide" sch_x=-95 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3106 N$6212 N$6211 "Straight Waveguide" sch_x=-95 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3107 N$6214 N$6213 "Straight Waveguide" sch_x=-95 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3108 N$6216 N$6215 "Straight Waveguide" sch_x=-95 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3109 N$6218 N$6217 "Straight Waveguide" sch_x=-95 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3110 N$6220 N$6219 "Straight Waveguide" sch_x=-95 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3111 N$6222 N$6221 "Straight Waveguide" sch_x=-95 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3112 N$6224 N$6223 "Straight Waveguide" sch_x=-95 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3113 N$6226 N$6225 "Straight Waveguide" sch_x=-95 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3114 N$6228 N$6227 "Straight Waveguide" sch_x=-95 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3115 N$6230 N$6229 "Straight Waveguide" sch_x=-95 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3116 N$6232 N$6231 "Straight Waveguide" sch_x=-95 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3117 N$6234 N$6233 "Straight Waveguide" sch_x=-95 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3118 N$6236 N$6235 "Straight Waveguide" sch_x=-95 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3119 N$6238 N$6237 "Straight Waveguide" sch_x=-95 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3120 N$6240 N$6239 "Straight Waveguide" sch_x=-95 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3121 N$6242 N$6241 "Straight Waveguide" sch_x=-93 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3122 N$6244 N$6243 "Straight Waveguide" sch_x=-93 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3123 N$6246 N$6245 "Straight Waveguide" sch_x=-93 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3124 N$6248 N$6247 "Straight Waveguide" sch_x=-93 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3125 N$6250 N$6249 "Straight Waveguide" sch_x=-93 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3126 N$6252 N$6251 "Straight Waveguide" sch_x=-93 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3127 N$6254 N$6253 "Straight Waveguide" sch_x=-93 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3128 N$6256 N$6255 "Straight Waveguide" sch_x=-93 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3129 N$6258 N$6257 "Straight Waveguide" sch_x=-93 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3130 N$6260 N$6259 "Straight Waveguide" sch_x=-93 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3131 N$6262 N$6261 "Straight Waveguide" sch_x=-93 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3132 N$6264 N$6263 "Straight Waveguide" sch_x=-93 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3133 N$6266 N$6265 "Straight Waveguide" sch_x=-93 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3134 N$6268 N$6267 "Straight Waveguide" sch_x=-93 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3135 N$6270 N$6269 "Straight Waveguide" sch_x=-93 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3136 N$6272 N$6271 "Straight Waveguide" sch_x=-93 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3137 N$6274 N$6273 "Straight Waveguide" sch_x=-93 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3138 N$6276 N$6275 "Straight Waveguide" sch_x=-93 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3139 N$6278 N$6277 "Straight Waveguide" sch_x=-93 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3140 N$6280 N$6279 "Straight Waveguide" sch_x=-93 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3141 N$6282 N$6281 "Straight Waveguide" sch_x=-93 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3142 N$6284 N$6283 "Straight Waveguide" sch_x=-93 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3143 N$6286 N$6285 "Straight Waveguide" sch_x=-93 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3144 N$6288 N$6287 "Straight Waveguide" sch_x=-93 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3145 N$6290 N$6289 "Straight Waveguide" sch_x=-93 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3146 N$6292 N$6291 "Straight Waveguide" sch_x=-93 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3147 N$6294 N$6293 "Straight Waveguide" sch_x=-93 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3148 N$6296 N$6295 "Straight Waveguide" sch_x=-93 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3149 N$6298 N$6297 "Straight Waveguide" sch_x=-93 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3150 N$6300 N$6299 "Straight Waveguide" sch_x=-93 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3151 N$6302 N$6301 "Straight Waveguide" sch_x=-91 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3152 N$6304 N$6303 "Straight Waveguide" sch_x=-91 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3153 N$6306 N$6305 "Straight Waveguide" sch_x=-91 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3154 N$6308 N$6307 "Straight Waveguide" sch_x=-91 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3155 N$6310 N$6309 "Straight Waveguide" sch_x=-91 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3156 N$6312 N$6311 "Straight Waveguide" sch_x=-91 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3157 N$6314 N$6313 "Straight Waveguide" sch_x=-91 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3158 N$6316 N$6315 "Straight Waveguide" sch_x=-91 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3159 N$6318 N$6317 "Straight Waveguide" sch_x=-91 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3160 N$6320 N$6319 "Straight Waveguide" sch_x=-91 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3161 N$6322 N$6321 "Straight Waveguide" sch_x=-91 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3162 N$6324 N$6323 "Straight Waveguide" sch_x=-91 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3163 N$6326 N$6325 "Straight Waveguide" sch_x=-91 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3164 N$6328 N$6327 "Straight Waveguide" sch_x=-91 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3165 N$6330 N$6329 "Straight Waveguide" sch_x=-91 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3166 N$6332 N$6331 "Straight Waveguide" sch_x=-91 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3167 N$6334 N$6333 "Straight Waveguide" sch_x=-91 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3168 N$6336 N$6335 "Straight Waveguide" sch_x=-91 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3169 N$6338 N$6337 "Straight Waveguide" sch_x=-91 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3170 N$6340 N$6339 "Straight Waveguide" sch_x=-91 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3171 N$6342 N$6341 "Straight Waveguide" sch_x=-91 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3172 N$6344 N$6343 "Straight Waveguide" sch_x=-91 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3173 N$6346 N$6345 "Straight Waveguide" sch_x=-91 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3174 N$6348 N$6347 "Straight Waveguide" sch_x=-91 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3175 N$6350 N$6349 "Straight Waveguide" sch_x=-91 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3176 N$6352 N$6351 "Straight Waveguide" sch_x=-91 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3177 N$6354 N$6353 "Straight Waveguide" sch_x=-91 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3178 N$6356 N$6355 "Straight Waveguide" sch_x=-91 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3179 N$6358 N$6357 "Straight Waveguide" sch_x=-89 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3180 N$6360 N$6359 "Straight Waveguide" sch_x=-89 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3181 N$6362 N$6361 "Straight Waveguide" sch_x=-89 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3182 N$6364 N$6363 "Straight Waveguide" sch_x=-89 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3183 N$6366 N$6365 "Straight Waveguide" sch_x=-89 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3184 N$6368 N$6367 "Straight Waveguide" sch_x=-89 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3185 N$6370 N$6369 "Straight Waveguide" sch_x=-89 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3186 N$6372 N$6371 "Straight Waveguide" sch_x=-89 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3187 N$6374 N$6373 "Straight Waveguide" sch_x=-89 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3188 N$6376 N$6375 "Straight Waveguide" sch_x=-89 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3189 N$6378 N$6377 "Straight Waveguide" sch_x=-89 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3190 N$6380 N$6379 "Straight Waveguide" sch_x=-89 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3191 N$6382 N$6381 "Straight Waveguide" sch_x=-89 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3192 N$6384 N$6383 "Straight Waveguide" sch_x=-89 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3193 N$6386 N$6385 "Straight Waveguide" sch_x=-89 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3194 N$6388 N$6387 "Straight Waveguide" sch_x=-89 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3195 N$6390 N$6389 "Straight Waveguide" sch_x=-89 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3196 N$6392 N$6391 "Straight Waveguide" sch_x=-89 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3197 N$6394 N$6393 "Straight Waveguide" sch_x=-89 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3198 N$6396 N$6395 "Straight Waveguide" sch_x=-89 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3199 N$6398 N$6397 "Straight Waveguide" sch_x=-89 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3200 N$6400 N$6399 "Straight Waveguide" sch_x=-89 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3201 N$6402 N$6401 "Straight Waveguide" sch_x=-89 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3202 N$6404 N$6403 "Straight Waveguide" sch_x=-89 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3203 N$6406 N$6405 "Straight Waveguide" sch_x=-89 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3204 N$6408 N$6407 "Straight Waveguide" sch_x=-89 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3205 N$6410 N$6409 "Straight Waveguide" sch_x=-87 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3206 N$6412 N$6411 "Straight Waveguide" sch_x=-87 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3207 N$6414 N$6413 "Straight Waveguide" sch_x=-87 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3208 N$6416 N$6415 "Straight Waveguide" sch_x=-87 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3209 N$6418 N$6417 "Straight Waveguide" sch_x=-87 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3210 N$6420 N$6419 "Straight Waveguide" sch_x=-87 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3211 N$6422 N$6421 "Straight Waveguide" sch_x=-87 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3212 N$6424 N$6423 "Straight Waveguide" sch_x=-87 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3213 N$6426 N$6425 "Straight Waveguide" sch_x=-87 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3214 N$6428 N$6427 "Straight Waveguide" sch_x=-87 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3215 N$6430 N$6429 "Straight Waveguide" sch_x=-87 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3216 N$6432 N$6431 "Straight Waveguide" sch_x=-87 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3217 N$6434 N$6433 "Straight Waveguide" sch_x=-87 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3218 N$6436 N$6435 "Straight Waveguide" sch_x=-87 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3219 N$6438 N$6437 "Straight Waveguide" sch_x=-87 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3220 N$6440 N$6439 "Straight Waveguide" sch_x=-87 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3221 N$6442 N$6441 "Straight Waveguide" sch_x=-87 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3222 N$6444 N$6443 "Straight Waveguide" sch_x=-87 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3223 N$6446 N$6445 "Straight Waveguide" sch_x=-87 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3224 N$6448 N$6447 "Straight Waveguide" sch_x=-87 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3225 N$6450 N$6449 "Straight Waveguide" sch_x=-87 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3226 N$6452 N$6451 "Straight Waveguide" sch_x=-87 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3227 N$6454 N$6453 "Straight Waveguide" sch_x=-87 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3228 N$6456 N$6455 "Straight Waveguide" sch_x=-87 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3229 N$6458 N$6457 "Straight Waveguide" sch_x=-85 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3230 N$6460 N$6459 "Straight Waveguide" sch_x=-85 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3231 N$6462 N$6461 "Straight Waveguide" sch_x=-85 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3232 N$6464 N$6463 "Straight Waveguide" sch_x=-85 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3233 N$6466 N$6465 "Straight Waveguide" sch_x=-85 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3234 N$6468 N$6467 "Straight Waveguide" sch_x=-85 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3235 N$6470 N$6469 "Straight Waveguide" sch_x=-85 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3236 N$6472 N$6471 "Straight Waveguide" sch_x=-85 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3237 N$6474 N$6473 "Straight Waveguide" sch_x=-85 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3238 N$6476 N$6475 "Straight Waveguide" sch_x=-85 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3239 N$6478 N$6477 "Straight Waveguide" sch_x=-85 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3240 N$6480 N$6479 "Straight Waveguide" sch_x=-85 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3241 N$6482 N$6481 "Straight Waveguide" sch_x=-85 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3242 N$6484 N$6483 "Straight Waveguide" sch_x=-85 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3243 N$6486 N$6485 "Straight Waveguide" sch_x=-85 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3244 N$6488 N$6487 "Straight Waveguide" sch_x=-85 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3245 N$6490 N$6489 "Straight Waveguide" sch_x=-85 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3246 N$6492 N$6491 "Straight Waveguide" sch_x=-85 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3247 N$6494 N$6493 "Straight Waveguide" sch_x=-85 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3248 N$6496 N$6495 "Straight Waveguide" sch_x=-85 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3249 N$6498 N$6497 "Straight Waveguide" sch_x=-85 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3250 N$6500 N$6499 "Straight Waveguide" sch_x=-85 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3251 N$6502 N$6501 "Straight Waveguide" sch_x=-83 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3252 N$6504 N$6503 "Straight Waveguide" sch_x=-83 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3253 N$6506 N$6505 "Straight Waveguide" sch_x=-83 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3254 N$6508 N$6507 "Straight Waveguide" sch_x=-83 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3255 N$6510 N$6509 "Straight Waveguide" sch_x=-83 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3256 N$6512 N$6511 "Straight Waveguide" sch_x=-83 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3257 N$6514 N$6513 "Straight Waveguide" sch_x=-83 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3258 N$6516 N$6515 "Straight Waveguide" sch_x=-83 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3259 N$6518 N$6517 "Straight Waveguide" sch_x=-83 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3260 N$6520 N$6519 "Straight Waveguide" sch_x=-83 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3261 N$6522 N$6521 "Straight Waveguide" sch_x=-83 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3262 N$6524 N$6523 "Straight Waveguide" sch_x=-83 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3263 N$6526 N$6525 "Straight Waveguide" sch_x=-83 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3264 N$6528 N$6527 "Straight Waveguide" sch_x=-83 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3265 N$6530 N$6529 "Straight Waveguide" sch_x=-83 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3266 N$6532 N$6531 "Straight Waveguide" sch_x=-83 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3267 N$6534 N$6533 "Straight Waveguide" sch_x=-83 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3268 N$6536 N$6535 "Straight Waveguide" sch_x=-83 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3269 N$6538 N$6537 "Straight Waveguide" sch_x=-83 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3270 N$6540 N$6539 "Straight Waveguide" sch_x=-83 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3271 N$6542 N$6541 "Straight Waveguide" sch_x=-81 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3272 N$6544 N$6543 "Straight Waveguide" sch_x=-81 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3273 N$6546 N$6545 "Straight Waveguide" sch_x=-81 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3274 N$6548 N$6547 "Straight Waveguide" sch_x=-81 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3275 N$6550 N$6549 "Straight Waveguide" sch_x=-81 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3276 N$6552 N$6551 "Straight Waveguide" sch_x=-81 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3277 N$6554 N$6553 "Straight Waveguide" sch_x=-81 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3278 N$6556 N$6555 "Straight Waveguide" sch_x=-81 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3279 N$6558 N$6557 "Straight Waveguide" sch_x=-81 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3280 N$6560 N$6559 "Straight Waveguide" sch_x=-81 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3281 N$6562 N$6561 "Straight Waveguide" sch_x=-81 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3282 N$6564 N$6563 "Straight Waveguide" sch_x=-81 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3283 N$6566 N$6565 "Straight Waveguide" sch_x=-81 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3284 N$6568 N$6567 "Straight Waveguide" sch_x=-81 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3285 N$6570 N$6569 "Straight Waveguide" sch_x=-81 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3286 N$6572 N$6571 "Straight Waveguide" sch_x=-81 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3287 N$6574 N$6573 "Straight Waveguide" sch_x=-81 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3288 N$6576 N$6575 "Straight Waveguide" sch_x=-81 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3289 N$6578 N$6577 "Straight Waveguide" sch_x=-79 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3290 N$6580 N$6579 "Straight Waveguide" sch_x=-79 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3291 N$6582 N$6581 "Straight Waveguide" sch_x=-79 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3292 N$6584 N$6583 "Straight Waveguide" sch_x=-79 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3293 N$6586 N$6585 "Straight Waveguide" sch_x=-79 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3294 N$6588 N$6587 "Straight Waveguide" sch_x=-79 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3295 N$6590 N$6589 "Straight Waveguide" sch_x=-79 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3296 N$6592 N$6591 "Straight Waveguide" sch_x=-79 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3297 N$6594 N$6593 "Straight Waveguide" sch_x=-79 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3298 N$6596 N$6595 "Straight Waveguide" sch_x=-79 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3299 N$6598 N$6597 "Straight Waveguide" sch_x=-79 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3300 N$6600 N$6599 "Straight Waveguide" sch_x=-79 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3301 N$6602 N$6601 "Straight Waveguide" sch_x=-79 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3302 N$6604 N$6603 "Straight Waveguide" sch_x=-79 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3303 N$6606 N$6605 "Straight Waveguide" sch_x=-79 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3304 N$6608 N$6607 "Straight Waveguide" sch_x=-79 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3305 N$6610 N$6609 "Straight Waveguide" sch_x=-77 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3306 N$6612 N$6611 "Straight Waveguide" sch_x=-77 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3307 N$6614 N$6613 "Straight Waveguide" sch_x=-77 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3308 N$6616 N$6615 "Straight Waveguide" sch_x=-77 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3309 N$6618 N$6617 "Straight Waveguide" sch_x=-77 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3310 N$6620 N$6619 "Straight Waveguide" sch_x=-77 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3311 N$6622 N$6621 "Straight Waveguide" sch_x=-77 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3312 N$6624 N$6623 "Straight Waveguide" sch_x=-77 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3313 N$6626 N$6625 "Straight Waveguide" sch_x=-77 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3314 N$6628 N$6627 "Straight Waveguide" sch_x=-77 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3315 N$6630 N$6629 "Straight Waveguide" sch_x=-77 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3316 N$6632 N$6631 "Straight Waveguide" sch_x=-77 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3317 N$6634 N$6633 "Straight Waveguide" sch_x=-77 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3318 N$6636 N$6635 "Straight Waveguide" sch_x=-77 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3319 N$6638 N$6637 "Straight Waveguide" sch_x=-75 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3320 N$6640 N$6639 "Straight Waveguide" sch_x=-75 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3321 N$6642 N$6641 "Straight Waveguide" sch_x=-75 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3322 N$6644 N$6643 "Straight Waveguide" sch_x=-75 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3323 N$6646 N$6645 "Straight Waveguide" sch_x=-75 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3324 N$6648 N$6647 "Straight Waveguide" sch_x=-75 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3325 N$6650 N$6649 "Straight Waveguide" sch_x=-75 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3326 N$6652 N$6651 "Straight Waveguide" sch_x=-75 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3327 N$6654 N$6653 "Straight Waveguide" sch_x=-75 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3328 N$6656 N$6655 "Straight Waveguide" sch_x=-75 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3329 N$6658 N$6657 "Straight Waveguide" sch_x=-75 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3330 N$6660 N$6659 "Straight Waveguide" sch_x=-75 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3331 N$6662 N$6661 "Straight Waveguide" sch_x=-73 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3332 N$6664 N$6663 "Straight Waveguide" sch_x=-73 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3333 N$6666 N$6665 "Straight Waveguide" sch_x=-73 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3334 N$6668 N$6667 "Straight Waveguide" sch_x=-73 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3335 N$6670 N$6669 "Straight Waveguide" sch_x=-73 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3336 N$6672 N$6671 "Straight Waveguide" sch_x=-73 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3337 N$6674 N$6673 "Straight Waveguide" sch_x=-73 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3338 N$6676 N$6675 "Straight Waveguide" sch_x=-73 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3339 N$6678 N$6677 "Straight Waveguide" sch_x=-73 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3340 N$6680 N$6679 "Straight Waveguide" sch_x=-73 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3341 N$6682 N$6681 "Straight Waveguide" sch_x=-71 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3342 N$6684 N$6683 "Straight Waveguide" sch_x=-71 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3343 N$6686 N$6685 "Straight Waveguide" sch_x=-71 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3344 N$6688 N$6687 "Straight Waveguide" sch_x=-71 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3345 N$6690 N$6689 "Straight Waveguide" sch_x=-71 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3346 N$6692 N$6691 "Straight Waveguide" sch_x=-71 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3347 N$6694 N$6693 "Straight Waveguide" sch_x=-71 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3348 N$6696 N$6695 "Straight Waveguide" sch_x=-71 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3349 N$6698 N$6697 "Straight Waveguide" sch_x=-69 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3350 N$6700 N$6699 "Straight Waveguide" sch_x=-69 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3351 N$6702 N$6701 "Straight Waveguide" sch_x=-69 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3352 N$6704 N$6703 "Straight Waveguide" sch_x=-69 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3353 N$6706 N$6705 "Straight Waveguide" sch_x=-69 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3354 N$6708 N$6707 "Straight Waveguide" sch_x=-69 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3355 N$6710 N$6709 "Straight Waveguide" sch_x=-67 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3356 N$6712 N$6711 "Straight Waveguide" sch_x=-67 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3357 N$6714 N$6713 "Straight Waveguide" sch_x=-67 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3358 N$6716 N$6715 "Straight Waveguide" sch_x=-67 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3359 N$6718 N$6717 "Straight Waveguide" sch_x=-65 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3360 N$6720 N$6719 "Straight Waveguide" sch_x=-65 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3361 N$6721 N$6722 "Straight Waveguide" sch_x=-93 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3362 N$6723 N$6724 "Straight Waveguide" sch_x=-92 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3363 N$6725 N$6726 "Straight Waveguide" sch_x=-91 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3364 N$6727 N$6728 "Straight Waveguide" sch_x=-90 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3365 N$6729 N$6730 "Straight Waveguide" sch_x=-89 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3366 N$6731 N$6732 "Straight Waveguide" sch_x=-88 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3367 N$6733 N$6734 "Straight Waveguide" sch_x=-87 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3368 N$6735 N$6736 "Straight Waveguide" sch_x=-86 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3369 N$6737 N$6738 "Straight Waveguide" sch_x=-85 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3370 N$6739 N$6740 "Straight Waveguide" sch_x=-84 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3371 N$6741 N$6742 "Straight Waveguide" sch_x=-83 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3372 N$6743 N$6744 "Straight Waveguide" sch_x=-82 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3373 N$6745 N$6746 "Straight Waveguide" sch_x=-81 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3374 N$6747 N$6748 "Straight Waveguide" sch_x=-80 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3375 N$6749 N$6750 "Straight Waveguide" sch_x=-79 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3376 N$6751 N$6752 "Straight Waveguide" sch_x=-78 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3377 N$6753 N$6754 "Straight Waveguide" sch_x=-77 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3378 N$6755 N$6756 "Straight Waveguide" sch_x=-76 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3379 N$6757 N$6758 "Straight Waveguide" sch_x=-75 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3380 N$6759 N$6760 "Straight Waveguide" sch_x=-74 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3381 N$6761 N$6762 "Straight Waveguide" sch_x=-73 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3382 N$6763 N$6764 "Straight Waveguide" sch_x=-72 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3383 N$6765 N$6766 "Straight Waveguide" sch_x=-71 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3384 N$6767 N$6768 "Straight Waveguide" sch_x=-70 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3385 N$6769 N$6770 "Straight Waveguide" sch_x=-69 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3386 N$6771 N$6772 "Straight Waveguide" sch_x=-68 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3387 N$6773 N$6774 "Straight Waveguide" sch_x=-67 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3388 N$6775 N$6776 "Straight Waveguide" sch_x=-66 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3389 N$6777 N$6778 "Straight Waveguide" sch_x=-65 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3390 N$6779 N$6780 "Straight Waveguide" sch_x=-64 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3391 N$6781 N$6782 "Straight Waveguide" sch_x=-63 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3392 N$6783 N$6784 "Straight Waveguide" sch_x=-63 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3393 N$6785 N$6786 "Straight Waveguide" sch_x=-64 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3394 N$6787 N$6788 "Straight Waveguide" sch_x=-65 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3395 N$6789 N$6790 "Straight Waveguide" sch_x=-66 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3396 N$6791 N$6792 "Straight Waveguide" sch_x=-67 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3397 N$6793 N$6794 "Straight Waveguide" sch_x=-68 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3398 N$6795 N$6796 "Straight Waveguide" sch_x=-69 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3399 N$6797 N$6798 "Straight Waveguide" sch_x=-70 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3400 N$6799 N$6800 "Straight Waveguide" sch_x=-71 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3401 N$6801 N$6802 "Straight Waveguide" sch_x=-72 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3402 N$6803 N$6804 "Straight Waveguide" sch_x=-73 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3403 N$6805 N$6806 "Straight Waveguide" sch_x=-74 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3404 N$6807 N$6808 "Straight Waveguide" sch_x=-75 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3405 N$6809 N$6810 "Straight Waveguide" sch_x=-76 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3406 N$6811 N$6812 "Straight Waveguide" sch_x=-77 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3407 N$6813 N$6814 "Straight Waveguide" sch_x=-78 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3408 N$6815 N$6816 "Straight Waveguide" sch_x=-79 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3409 N$6817 N$6818 "Straight Waveguide" sch_x=-80 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3410 N$6819 N$6820 "Straight Waveguide" sch_x=-81 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3411 N$6821 N$6822 "Straight Waveguide" sch_x=-82 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3412 N$6823 N$6824 "Straight Waveguide" sch_x=-83 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3413 N$6825 N$6826 "Straight Waveguide" sch_x=-84 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3414 N$6827 N$6828 "Straight Waveguide" sch_x=-85 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3415 N$6829 N$6830 "Straight Waveguide" sch_x=-86 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3416 N$6831 N$6832 "Straight Waveguide" sch_x=-87 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3417 N$6833 N$6834 "Straight Waveguide" sch_x=-88 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3418 N$6835 N$6836 "Straight Waveguide" sch_x=-89 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3419 N$6837 N$6838 "Straight Waveguide" sch_x=-90 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3420 N$6839 N$6840 "Straight Waveguide" sch_x=-91 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3421 N$6841 N$6842 "Straight Waveguide" sch_x=-92 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3422 N$6843 N$6844 "Straight Waveguide" sch_x=-93 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3423 N$6845 N$6846 "Straight Waveguide" sch_x=-94 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3424 N$6847 N$6848 "Straight Waveguide" sch_x=-94 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3425 N$6849 N$6850 "Straight Waveguide" sch_x=125 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3426 N$6851 N$6852 "Straight Waveguide" sch_x=125 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3427 N$6853 N$6854 "Straight Waveguide" sch_x=125 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3428 N$6855 N$6856 "Straight Waveguide" sch_x=125 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3429 N$6857 N$6858 "Straight Waveguide" sch_x=125 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3430 N$6859 N$6860 "Straight Waveguide" sch_x=125 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3431 N$6861 N$6862 "Straight Waveguide" sch_x=125 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3432 N$6863 N$6864 "Straight Waveguide" sch_x=125 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3433 N$6865 N$6866 "Straight Waveguide" sch_x=125 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3434 N$6867 N$6868 "Straight Waveguide" sch_x=125 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3435 N$6869 N$6870 "Straight Waveguide" sch_x=125 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3436 N$6871 N$6872 "Straight Waveguide" sch_x=125 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3437 N$6873 N$6874 "Straight Waveguide" sch_x=125 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3438 N$6875 N$6876 "Straight Waveguide" sch_x=125 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3439 N$6877 N$6878 "Straight Waveguide" sch_x=125 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3440 N$6879 N$6880 "Straight Waveguide" sch_x=125 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3441 N$6881 N$6882 "Straight Waveguide" sch_x=125 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3442 N$6883 N$6884 "Straight Waveguide" sch_x=125 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3443 N$6885 N$6886 "Straight Waveguide" sch_x=125 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3444 N$6887 N$6888 "Straight Waveguide" sch_x=125 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3445 N$6889 N$6890 "Straight Waveguide" sch_x=125 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3446 N$6891 N$6892 "Straight Waveguide" sch_x=125 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3447 N$6893 N$6894 "Straight Waveguide" sch_x=125 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3448 N$6895 N$6896 "Straight Waveguide" sch_x=125 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3449 N$6897 N$6898 "Straight Waveguide" sch_x=125 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3450 N$6899 N$6900 "Straight Waveguide" sch_x=125 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3451 N$6901 N$6902 "Straight Waveguide" sch_x=125 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3452 N$6903 N$6904 "Straight Waveguide" sch_x=125 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3453 N$6905 N$6906 "Straight Waveguide" sch_x=125 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3454 N$6907 N$6908 "Straight Waveguide" sch_x=125 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3455 N$6909 N$6910 "Straight Waveguide" sch_x=125 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3456 N$6911 N$6912 "Straight Waveguide" sch_x=125 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3457 N$6913 N$6914 "Straight Waveguide" sch_x=125 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3458 N$6915 N$6916 "Straight Waveguide" sch_x=125 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3459 N$6917 N$6918 "Straight Waveguide" sch_x=125 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3460 N$6919 N$6920 "Straight Waveguide" sch_x=125 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3461 N$6921 N$6922 "Straight Waveguide" sch_x=125 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3462 N$6923 N$6924 "Straight Waveguide" sch_x=125 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3463 N$6925 N$6926 "Straight Waveguide" sch_x=125 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3464 N$6927 N$6928 "Straight Waveguide" sch_x=125 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3465 N$6929 N$6930 "Straight Waveguide" sch_x=125 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3466 N$6931 N$6932 "Straight Waveguide" sch_x=125 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3467 N$6933 N$6934 "Straight Waveguide" sch_x=125 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3468 N$6935 N$6936 "Straight Waveguide" sch_x=125 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3469 N$6937 N$6938 "Straight Waveguide" sch_x=125 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3470 N$6939 N$6940 "Straight Waveguide" sch_x=125 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3471 N$6941 N$6942 "Straight Waveguide" sch_x=125 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3472 N$6943 N$6944 "Straight Waveguide" sch_x=125 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3473 N$6945 N$6946 "Straight Waveguide" sch_x=125 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3474 N$6947 N$6948 "Straight Waveguide" sch_x=125 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3475 N$6949 N$6950 "Straight Waveguide" sch_x=125 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3476 N$6951 N$6952 "Straight Waveguide" sch_x=125 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3477 N$6953 N$6954 "Straight Waveguide" sch_x=125 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3478 N$6955 N$6956 "Straight Waveguide" sch_x=125 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3479 N$6957 N$6958 "Straight Waveguide" sch_x=125 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3480 N$6959 N$6960 "Straight Waveguide" sch_x=125 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3481 N$6961 N$6962 "Straight Waveguide" sch_x=125 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3482 N$6963 N$6964 "Straight Waveguide" sch_x=125 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3483 N$6965 N$6966 "Straight Waveguide" sch_x=125 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3484 N$6967 N$6968 "Straight Waveguide" sch_x=125 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3485 N$6969 N$6970 "Straight Waveguide" sch_x=125 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3486 N$6971 N$6972 "Straight Waveguide" sch_x=125 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3487 N$6973 N$6974 "Straight Waveguide" sch_x=123 sch_y=29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3488 N$6975 N$6976 "Straight Waveguide" sch_x=123 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3489 N$6977 N$6978 "Straight Waveguide" sch_x=123 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3490 N$6979 N$6980 "Straight Waveguide" sch_x=123 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3491 N$6981 N$6982 "Straight Waveguide" sch_x=123 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3492 N$6983 N$6984 "Straight Waveguide" sch_x=123 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3493 N$6985 N$6986 "Straight Waveguide" sch_x=123 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3494 N$6987 N$6988 "Straight Waveguide" sch_x=123 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3495 N$6989 N$6990 "Straight Waveguide" sch_x=123 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3496 N$6991 N$6992 "Straight Waveguide" sch_x=123 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3497 N$6993 N$6994 "Straight Waveguide" sch_x=123 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3498 N$6995 N$6996 "Straight Waveguide" sch_x=123 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3499 N$6997 N$6998 "Straight Waveguide" sch_x=123 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3500 N$6999 N$7000 "Straight Waveguide" sch_x=123 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3501 N$7001 N$7002 "Straight Waveguide" sch_x=123 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3502 N$7003 N$7004 "Straight Waveguide" sch_x=123 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3503 N$7005 N$7006 "Straight Waveguide" sch_x=123 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3504 N$7007 N$7008 "Straight Waveguide" sch_x=123 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3505 N$7009 N$7010 "Straight Waveguide" sch_x=123 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3506 N$7011 N$7012 "Straight Waveguide" sch_x=123 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3507 N$7013 N$7014 "Straight Waveguide" sch_x=123 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3508 N$7015 N$7016 "Straight Waveguide" sch_x=123 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3509 N$7017 N$7018 "Straight Waveguide" sch_x=123 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3510 N$7019 N$7020 "Straight Waveguide" sch_x=123 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3511 N$7021 N$7022 "Straight Waveguide" sch_x=123 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3512 N$7023 N$7024 "Straight Waveguide" sch_x=123 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3513 N$7025 N$7026 "Straight Waveguide" sch_x=123 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3514 N$7027 N$7028 "Straight Waveguide" sch_x=123 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3515 N$7029 N$7030 "Straight Waveguide" sch_x=123 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3516 N$7031 N$7032 "Straight Waveguide" sch_x=123 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3517 N$7033 N$7034 "Straight Waveguide" sch_x=123 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3518 N$7035 N$7036 "Straight Waveguide" sch_x=123 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3519 N$7037 N$7038 "Straight Waveguide" sch_x=123 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3520 N$7039 N$7040 "Straight Waveguide" sch_x=123 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3521 N$7041 N$7042 "Straight Waveguide" sch_x=123 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3522 N$7043 N$7044 "Straight Waveguide" sch_x=123 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3523 N$7045 N$7046 "Straight Waveguide" sch_x=123 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3524 N$7047 N$7048 "Straight Waveguide" sch_x=123 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3525 N$7049 N$7050 "Straight Waveguide" sch_x=123 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3526 N$7051 N$7052 "Straight Waveguide" sch_x=123 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3527 N$7053 N$7054 "Straight Waveguide" sch_x=123 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3528 N$7055 N$7056 "Straight Waveguide" sch_x=123 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3529 N$7057 N$7058 "Straight Waveguide" sch_x=123 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3530 N$7059 N$7060 "Straight Waveguide" sch_x=123 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3531 N$7061 N$7062 "Straight Waveguide" sch_x=123 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3532 N$7063 N$7064 "Straight Waveguide" sch_x=123 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3533 N$7065 N$7066 "Straight Waveguide" sch_x=123 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3534 N$7067 N$7068 "Straight Waveguide" sch_x=123 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3535 N$7069 N$7070 "Straight Waveguide" sch_x=123 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3536 N$7071 N$7072 "Straight Waveguide" sch_x=123 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3537 N$7073 N$7074 "Straight Waveguide" sch_x=123 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3538 N$7075 N$7076 "Straight Waveguide" sch_x=123 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3539 N$7077 N$7078 "Straight Waveguide" sch_x=123 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3540 N$7079 N$7080 "Straight Waveguide" sch_x=123 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3541 N$7081 N$7082 "Straight Waveguide" sch_x=123 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3542 N$7083 N$7084 "Straight Waveguide" sch_x=123 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3543 N$7085 N$7086 "Straight Waveguide" sch_x=123 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3544 N$7087 N$7088 "Straight Waveguide" sch_x=123 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3545 N$7089 N$7090 "Straight Waveguide" sch_x=123 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3546 N$7091 N$7092 "Straight Waveguide" sch_x=123 sch_y=-29.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3547 N$7093 N$7094 "Straight Waveguide" sch_x=121 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3548 N$7095 N$7096 "Straight Waveguide" sch_x=121 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3549 N$7097 N$7098 "Straight Waveguide" sch_x=121 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3550 N$7099 N$7100 "Straight Waveguide" sch_x=121 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3551 N$7101 N$7102 "Straight Waveguide" sch_x=121 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3552 N$7103 N$7104 "Straight Waveguide" sch_x=121 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3553 N$7105 N$7106 "Straight Waveguide" sch_x=121 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3554 N$7107 N$7108 "Straight Waveguide" sch_x=121 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3555 N$7109 N$7110 "Straight Waveguide" sch_x=121 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3556 N$7111 N$7112 "Straight Waveguide" sch_x=121 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3557 N$7113 N$7114 "Straight Waveguide" sch_x=121 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3558 N$7115 N$7116 "Straight Waveguide" sch_x=121 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3559 N$7117 N$7118 "Straight Waveguide" sch_x=121 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3560 N$7119 N$7120 "Straight Waveguide" sch_x=121 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3561 N$7121 N$7122 "Straight Waveguide" sch_x=121 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3562 N$7123 N$7124 "Straight Waveguide" sch_x=121 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3563 N$7125 N$7126 "Straight Waveguide" sch_x=121 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3564 N$7127 N$7128 "Straight Waveguide" sch_x=121 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3565 N$7129 N$7130 "Straight Waveguide" sch_x=121 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3566 N$7131 N$7132 "Straight Waveguide" sch_x=121 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3567 N$7133 N$7134 "Straight Waveguide" sch_x=121 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3568 N$7135 N$7136 "Straight Waveguide" sch_x=121 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3569 N$7137 N$7138 "Straight Waveguide" sch_x=121 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3570 N$7139 N$7140 "Straight Waveguide" sch_x=121 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3571 N$7141 N$7142 "Straight Waveguide" sch_x=121 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3572 N$7143 N$7144 "Straight Waveguide" sch_x=121 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3573 N$7145 N$7146 "Straight Waveguide" sch_x=121 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3574 N$7147 N$7148 "Straight Waveguide" sch_x=121 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3575 N$7149 N$7150 "Straight Waveguide" sch_x=121 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3576 N$7151 N$7152 "Straight Waveguide" sch_x=121 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3577 N$7153 N$7154 "Straight Waveguide" sch_x=121 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3578 N$7155 N$7156 "Straight Waveguide" sch_x=121 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3579 N$7157 N$7158 "Straight Waveguide" sch_x=121 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3580 N$7159 N$7160 "Straight Waveguide" sch_x=121 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3581 N$7161 N$7162 "Straight Waveguide" sch_x=121 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3582 N$7163 N$7164 "Straight Waveguide" sch_x=121 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3583 N$7165 N$7166 "Straight Waveguide" sch_x=121 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3584 N$7167 N$7168 "Straight Waveguide" sch_x=121 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3585 N$7169 N$7170 "Straight Waveguide" sch_x=121 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3586 N$7171 N$7172 "Straight Waveguide" sch_x=121 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3587 N$7173 N$7174 "Straight Waveguide" sch_x=121 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3588 N$7175 N$7176 "Straight Waveguide" sch_x=121 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3589 N$7177 N$7178 "Straight Waveguide" sch_x=121 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3590 N$7179 N$7180 "Straight Waveguide" sch_x=121 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3591 N$7181 N$7182 "Straight Waveguide" sch_x=121 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3592 N$7183 N$7184 "Straight Waveguide" sch_x=121 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3593 N$7185 N$7186 "Straight Waveguide" sch_x=121 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3594 N$7187 N$7188 "Straight Waveguide" sch_x=121 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3595 N$7189 N$7190 "Straight Waveguide" sch_x=121 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3596 N$7191 N$7192 "Straight Waveguide" sch_x=121 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3597 N$7193 N$7194 "Straight Waveguide" sch_x=121 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3598 N$7195 N$7196 "Straight Waveguide" sch_x=121 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3599 N$7197 N$7198 "Straight Waveguide" sch_x=121 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3600 N$7199 N$7200 "Straight Waveguide" sch_x=121 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3601 N$7201 N$7202 "Straight Waveguide" sch_x=121 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3602 N$7203 N$7204 "Straight Waveguide" sch_x=121 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3603 N$7205 N$7206 "Straight Waveguide" sch_x=121 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3604 N$7207 N$7208 "Straight Waveguide" sch_x=121 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3605 N$7209 N$7210 "Straight Waveguide" sch_x=119 sch_y=27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3606 N$7211 N$7212 "Straight Waveguide" sch_x=119 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3607 N$7213 N$7214 "Straight Waveguide" sch_x=119 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3608 N$7215 N$7216 "Straight Waveguide" sch_x=119 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3609 N$7217 N$7218 "Straight Waveguide" sch_x=119 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3610 N$7219 N$7220 "Straight Waveguide" sch_x=119 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3611 N$7221 N$7222 "Straight Waveguide" sch_x=119 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3612 N$7223 N$7224 "Straight Waveguide" sch_x=119 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3613 N$7225 N$7226 "Straight Waveguide" sch_x=119 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3614 N$7227 N$7228 "Straight Waveguide" sch_x=119 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3615 N$7229 N$7230 "Straight Waveguide" sch_x=119 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3616 N$7231 N$7232 "Straight Waveguide" sch_x=119 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3617 N$7233 N$7234 "Straight Waveguide" sch_x=119 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3618 N$7235 N$7236 "Straight Waveguide" sch_x=119 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3619 N$7237 N$7238 "Straight Waveguide" sch_x=119 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3620 N$7239 N$7240 "Straight Waveguide" sch_x=119 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3621 N$7241 N$7242 "Straight Waveguide" sch_x=119 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3622 N$7243 N$7244 "Straight Waveguide" sch_x=119 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3623 N$7245 N$7246 "Straight Waveguide" sch_x=119 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3624 N$7247 N$7248 "Straight Waveguide" sch_x=119 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3625 N$7249 N$7250 "Straight Waveguide" sch_x=119 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3626 N$7251 N$7252 "Straight Waveguide" sch_x=119 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3627 N$7253 N$7254 "Straight Waveguide" sch_x=119 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3628 N$7255 N$7256 "Straight Waveguide" sch_x=119 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3629 N$7257 N$7258 "Straight Waveguide" sch_x=119 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3630 N$7259 N$7260 "Straight Waveguide" sch_x=119 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3631 N$7261 N$7262 "Straight Waveguide" sch_x=119 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3632 N$7263 N$7264 "Straight Waveguide" sch_x=119 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3633 N$7265 N$7266 "Straight Waveguide" sch_x=119 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3634 N$7267 N$7268 "Straight Waveguide" sch_x=119 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3635 N$7269 N$7270 "Straight Waveguide" sch_x=119 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3636 N$7271 N$7272 "Straight Waveguide" sch_x=119 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3637 N$7273 N$7274 "Straight Waveguide" sch_x=119 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3638 N$7275 N$7276 "Straight Waveguide" sch_x=119 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3639 N$7277 N$7278 "Straight Waveguide" sch_x=119 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3640 N$7279 N$7280 "Straight Waveguide" sch_x=119 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3641 N$7281 N$7282 "Straight Waveguide" sch_x=119 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3642 N$7283 N$7284 "Straight Waveguide" sch_x=119 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3643 N$7285 N$7286 "Straight Waveguide" sch_x=119 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3644 N$7287 N$7288 "Straight Waveguide" sch_x=119 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3645 N$7289 N$7290 "Straight Waveguide" sch_x=119 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3646 N$7291 N$7292 "Straight Waveguide" sch_x=119 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3647 N$7293 N$7294 "Straight Waveguide" sch_x=119 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3648 N$7295 N$7296 "Straight Waveguide" sch_x=119 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3649 N$7297 N$7298 "Straight Waveguide" sch_x=119 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3650 N$7299 N$7300 "Straight Waveguide" sch_x=119 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3651 N$7301 N$7302 "Straight Waveguide" sch_x=119 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3652 N$7303 N$7304 "Straight Waveguide" sch_x=119 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3653 N$7305 N$7306 "Straight Waveguide" sch_x=119 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3654 N$7307 N$7308 "Straight Waveguide" sch_x=119 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3655 N$7309 N$7310 "Straight Waveguide" sch_x=119 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3656 N$7311 N$7312 "Straight Waveguide" sch_x=119 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3657 N$7313 N$7314 "Straight Waveguide" sch_x=119 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3658 N$7315 N$7316 "Straight Waveguide" sch_x=119 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3659 N$7317 N$7318 "Straight Waveguide" sch_x=119 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3660 N$7319 N$7320 "Straight Waveguide" sch_x=119 sch_y=-27.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3661 N$7321 N$7322 "Straight Waveguide" sch_x=117 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3662 N$7323 N$7324 "Straight Waveguide" sch_x=117 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3663 N$7325 N$7326 "Straight Waveguide" sch_x=117 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3664 N$7327 N$7328 "Straight Waveguide" sch_x=117 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3665 N$7329 N$7330 "Straight Waveguide" sch_x=117 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3666 N$7331 N$7332 "Straight Waveguide" sch_x=117 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3667 N$7333 N$7334 "Straight Waveguide" sch_x=117 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3668 N$7335 N$7336 "Straight Waveguide" sch_x=117 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3669 N$7337 N$7338 "Straight Waveguide" sch_x=117 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3670 N$7339 N$7340 "Straight Waveguide" sch_x=117 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3671 N$7341 N$7342 "Straight Waveguide" sch_x=117 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3672 N$7343 N$7344 "Straight Waveguide" sch_x=117 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3673 N$7345 N$7346 "Straight Waveguide" sch_x=117 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3674 N$7347 N$7348 "Straight Waveguide" sch_x=117 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3675 N$7349 N$7350 "Straight Waveguide" sch_x=117 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3676 N$7351 N$7352 "Straight Waveguide" sch_x=117 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3677 N$7353 N$7354 "Straight Waveguide" sch_x=117 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3678 N$7355 N$7356 "Straight Waveguide" sch_x=117 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3679 N$7357 N$7358 "Straight Waveguide" sch_x=117 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3680 N$7359 N$7360 "Straight Waveguide" sch_x=117 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3681 N$7361 N$7362 "Straight Waveguide" sch_x=117 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3682 N$7363 N$7364 "Straight Waveguide" sch_x=117 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3683 N$7365 N$7366 "Straight Waveguide" sch_x=117 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3684 N$7367 N$7368 "Straight Waveguide" sch_x=117 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3685 N$7369 N$7370 "Straight Waveguide" sch_x=117 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3686 N$7371 N$7372 "Straight Waveguide" sch_x=117 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3687 N$7373 N$7374 "Straight Waveguide" sch_x=117 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3688 N$7375 N$7376 "Straight Waveguide" sch_x=117 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3689 N$7377 N$7378 "Straight Waveguide" sch_x=117 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3690 N$7379 N$7380 "Straight Waveguide" sch_x=117 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3691 N$7381 N$7382 "Straight Waveguide" sch_x=117 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3692 N$7383 N$7384 "Straight Waveguide" sch_x=117 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3693 N$7385 N$7386 "Straight Waveguide" sch_x=117 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3694 N$7387 N$7388 "Straight Waveguide" sch_x=117 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3695 N$7389 N$7390 "Straight Waveguide" sch_x=117 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3696 N$7391 N$7392 "Straight Waveguide" sch_x=117 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3697 N$7393 N$7394 "Straight Waveguide" sch_x=117 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3698 N$7395 N$7396 "Straight Waveguide" sch_x=117 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3699 N$7397 N$7398 "Straight Waveguide" sch_x=117 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3700 N$7399 N$7400 "Straight Waveguide" sch_x=117 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3701 N$7401 N$7402 "Straight Waveguide" sch_x=117 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3702 N$7403 N$7404 "Straight Waveguide" sch_x=117 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3703 N$7405 N$7406 "Straight Waveguide" sch_x=117 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3704 N$7407 N$7408 "Straight Waveguide" sch_x=117 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3705 N$7409 N$7410 "Straight Waveguide" sch_x=117 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3706 N$7411 N$7412 "Straight Waveguide" sch_x=117 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3707 N$7413 N$7414 "Straight Waveguide" sch_x=117 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3708 N$7415 N$7416 "Straight Waveguide" sch_x=117 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3709 N$7417 N$7418 "Straight Waveguide" sch_x=117 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3710 N$7419 N$7420 "Straight Waveguide" sch_x=117 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3711 N$7421 N$7422 "Straight Waveguide" sch_x=117 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3712 N$7423 N$7424 "Straight Waveguide" sch_x=117 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3713 N$7425 N$7426 "Straight Waveguide" sch_x=117 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3714 N$7427 N$7428 "Straight Waveguide" sch_x=117 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3715 N$7429 N$7430 "Straight Waveguide" sch_x=115 sch_y=25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3716 N$7431 N$7432 "Straight Waveguide" sch_x=115 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3717 N$7433 N$7434 "Straight Waveguide" sch_x=115 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3718 N$7435 N$7436 "Straight Waveguide" sch_x=115 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3719 N$7437 N$7438 "Straight Waveguide" sch_x=115 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3720 N$7439 N$7440 "Straight Waveguide" sch_x=115 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3721 N$7441 N$7442 "Straight Waveguide" sch_x=115 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3722 N$7443 N$7444 "Straight Waveguide" sch_x=115 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3723 N$7445 N$7446 "Straight Waveguide" sch_x=115 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3724 N$7447 N$7448 "Straight Waveguide" sch_x=115 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3725 N$7449 N$7450 "Straight Waveguide" sch_x=115 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3726 N$7451 N$7452 "Straight Waveguide" sch_x=115 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3727 N$7453 N$7454 "Straight Waveguide" sch_x=115 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3728 N$7455 N$7456 "Straight Waveguide" sch_x=115 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3729 N$7457 N$7458 "Straight Waveguide" sch_x=115 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3730 N$7459 N$7460 "Straight Waveguide" sch_x=115 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3731 N$7461 N$7462 "Straight Waveguide" sch_x=115 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3732 N$7463 N$7464 "Straight Waveguide" sch_x=115 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3733 N$7465 N$7466 "Straight Waveguide" sch_x=115 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3734 N$7467 N$7468 "Straight Waveguide" sch_x=115 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3735 N$7469 N$7470 "Straight Waveguide" sch_x=115 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3736 N$7471 N$7472 "Straight Waveguide" sch_x=115 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3737 N$7473 N$7474 "Straight Waveguide" sch_x=115 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3738 N$7475 N$7476 "Straight Waveguide" sch_x=115 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3739 N$7477 N$7478 "Straight Waveguide" sch_x=115 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3740 N$7479 N$7480 "Straight Waveguide" sch_x=115 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3741 N$7481 N$7482 "Straight Waveguide" sch_x=115 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3742 N$7483 N$7484 "Straight Waveguide" sch_x=115 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3743 N$7485 N$7486 "Straight Waveguide" sch_x=115 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3744 N$7487 N$7488 "Straight Waveguide" sch_x=115 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3745 N$7489 N$7490 "Straight Waveguide" sch_x=115 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3746 N$7491 N$7492 "Straight Waveguide" sch_x=115 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3747 N$7493 N$7494 "Straight Waveguide" sch_x=115 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3748 N$7495 N$7496 "Straight Waveguide" sch_x=115 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3749 N$7497 N$7498 "Straight Waveguide" sch_x=115 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3750 N$7499 N$7500 "Straight Waveguide" sch_x=115 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3751 N$7501 N$7502 "Straight Waveguide" sch_x=115 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3752 N$7503 N$7504 "Straight Waveguide" sch_x=115 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3753 N$7505 N$7506 "Straight Waveguide" sch_x=115 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3754 N$7507 N$7508 "Straight Waveguide" sch_x=115 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3755 N$7509 N$7510 "Straight Waveguide" sch_x=115 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3756 N$7511 N$7512 "Straight Waveguide" sch_x=115 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3757 N$7513 N$7514 "Straight Waveguide" sch_x=115 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3758 N$7515 N$7516 "Straight Waveguide" sch_x=115 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3759 N$7517 N$7518 "Straight Waveguide" sch_x=115 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3760 N$7519 N$7520 "Straight Waveguide" sch_x=115 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3761 N$7521 N$7522 "Straight Waveguide" sch_x=115 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3762 N$7523 N$7524 "Straight Waveguide" sch_x=115 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3763 N$7525 N$7526 "Straight Waveguide" sch_x=115 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3764 N$7527 N$7528 "Straight Waveguide" sch_x=115 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3765 N$7529 N$7530 "Straight Waveguide" sch_x=115 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3766 N$7531 N$7532 "Straight Waveguide" sch_x=115 sch_y=-25.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3767 N$7533 N$7534 "Straight Waveguide" sch_x=113 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3768 N$7535 N$7536 "Straight Waveguide" sch_x=113 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3769 N$7537 N$7538 "Straight Waveguide" sch_x=113 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3770 N$7539 N$7540 "Straight Waveguide" sch_x=113 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3771 N$7541 N$7542 "Straight Waveguide" sch_x=113 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3772 N$7543 N$7544 "Straight Waveguide" sch_x=113 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3773 N$7545 N$7546 "Straight Waveguide" sch_x=113 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3774 N$7547 N$7548 "Straight Waveguide" sch_x=113 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3775 N$7549 N$7550 "Straight Waveguide" sch_x=113 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3776 N$7551 N$7552 "Straight Waveguide" sch_x=113 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3777 N$7553 N$7554 "Straight Waveguide" sch_x=113 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3778 N$7555 N$7556 "Straight Waveguide" sch_x=113 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3779 N$7557 N$7558 "Straight Waveguide" sch_x=113 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3780 N$7559 N$7560 "Straight Waveguide" sch_x=113 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3781 N$7561 N$7562 "Straight Waveguide" sch_x=113 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3782 N$7563 N$7564 "Straight Waveguide" sch_x=113 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3783 N$7565 N$7566 "Straight Waveguide" sch_x=113 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3784 N$7567 N$7568 "Straight Waveguide" sch_x=113 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3785 N$7569 N$7570 "Straight Waveguide" sch_x=113 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3786 N$7571 N$7572 "Straight Waveguide" sch_x=113 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3787 N$7573 N$7574 "Straight Waveguide" sch_x=113 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3788 N$7575 N$7576 "Straight Waveguide" sch_x=113 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3789 N$7577 N$7578 "Straight Waveguide" sch_x=113 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3790 N$7579 N$7580 "Straight Waveguide" sch_x=113 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3791 N$7581 N$7582 "Straight Waveguide" sch_x=113 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3792 N$7583 N$7584 "Straight Waveguide" sch_x=113 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3793 N$7585 N$7586 "Straight Waveguide" sch_x=113 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3794 N$7587 N$7588 "Straight Waveguide" sch_x=113 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3795 N$7589 N$7590 "Straight Waveguide" sch_x=113 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3796 N$7591 N$7592 "Straight Waveguide" sch_x=113 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3797 N$7593 N$7594 "Straight Waveguide" sch_x=113 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3798 N$7595 N$7596 "Straight Waveguide" sch_x=113 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3799 N$7597 N$7598 "Straight Waveguide" sch_x=113 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3800 N$7599 N$7600 "Straight Waveguide" sch_x=113 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3801 N$7601 N$7602 "Straight Waveguide" sch_x=113 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3802 N$7603 N$7604 "Straight Waveguide" sch_x=113 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3803 N$7605 N$7606 "Straight Waveguide" sch_x=113 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3804 N$7607 N$7608 "Straight Waveguide" sch_x=113 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3805 N$7609 N$7610 "Straight Waveguide" sch_x=113 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3806 N$7611 N$7612 "Straight Waveguide" sch_x=113 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3807 N$7613 N$7614 "Straight Waveguide" sch_x=113 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3808 N$7615 N$7616 "Straight Waveguide" sch_x=113 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3809 N$7617 N$7618 "Straight Waveguide" sch_x=113 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3810 N$7619 N$7620 "Straight Waveguide" sch_x=113 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3811 N$7621 N$7622 "Straight Waveguide" sch_x=113 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3812 N$7623 N$7624 "Straight Waveguide" sch_x=113 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3813 N$7625 N$7626 "Straight Waveguide" sch_x=113 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3814 N$7627 N$7628 "Straight Waveguide" sch_x=113 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3815 N$7629 N$7630 "Straight Waveguide" sch_x=113 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3816 N$7631 N$7632 "Straight Waveguide" sch_x=113 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3817 N$7633 N$7634 "Straight Waveguide" sch_x=111 sch_y=23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3818 N$7635 N$7636 "Straight Waveguide" sch_x=111 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3819 N$7637 N$7638 "Straight Waveguide" sch_x=111 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3820 N$7639 N$7640 "Straight Waveguide" sch_x=111 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3821 N$7641 N$7642 "Straight Waveguide" sch_x=111 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3822 N$7643 N$7644 "Straight Waveguide" sch_x=111 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3823 N$7645 N$7646 "Straight Waveguide" sch_x=111 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3824 N$7647 N$7648 "Straight Waveguide" sch_x=111 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3825 N$7649 N$7650 "Straight Waveguide" sch_x=111 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3826 N$7651 N$7652 "Straight Waveguide" sch_x=111 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3827 N$7653 N$7654 "Straight Waveguide" sch_x=111 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3828 N$7655 N$7656 "Straight Waveguide" sch_x=111 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3829 N$7657 N$7658 "Straight Waveguide" sch_x=111 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3830 N$7659 N$7660 "Straight Waveguide" sch_x=111 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3831 N$7661 N$7662 "Straight Waveguide" sch_x=111 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3832 N$7663 N$7664 "Straight Waveguide" sch_x=111 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3833 N$7665 N$7666 "Straight Waveguide" sch_x=111 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3834 N$7667 N$7668 "Straight Waveguide" sch_x=111 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3835 N$7669 N$7670 "Straight Waveguide" sch_x=111 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3836 N$7671 N$7672 "Straight Waveguide" sch_x=111 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3837 N$7673 N$7674 "Straight Waveguide" sch_x=111 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3838 N$7675 N$7676 "Straight Waveguide" sch_x=111 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3839 N$7677 N$7678 "Straight Waveguide" sch_x=111 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3840 N$7679 N$7680 "Straight Waveguide" sch_x=111 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3841 N$7681 N$7682 "Straight Waveguide" sch_x=111 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3842 N$7683 N$7684 "Straight Waveguide" sch_x=111 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3843 N$7685 N$7686 "Straight Waveguide" sch_x=111 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3844 N$7687 N$7688 "Straight Waveguide" sch_x=111 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3845 N$7689 N$7690 "Straight Waveguide" sch_x=111 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3846 N$7691 N$7692 "Straight Waveguide" sch_x=111 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3847 N$7693 N$7694 "Straight Waveguide" sch_x=111 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3848 N$7695 N$7696 "Straight Waveguide" sch_x=111 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3849 N$7697 N$7698 "Straight Waveguide" sch_x=111 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3850 N$7699 N$7700 "Straight Waveguide" sch_x=111 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3851 N$7701 N$7702 "Straight Waveguide" sch_x=111 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3852 N$7703 N$7704 "Straight Waveguide" sch_x=111 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3853 N$7705 N$7706 "Straight Waveguide" sch_x=111 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3854 N$7707 N$7708 "Straight Waveguide" sch_x=111 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3855 N$7709 N$7710 "Straight Waveguide" sch_x=111 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3856 N$7711 N$7712 "Straight Waveguide" sch_x=111 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3857 N$7713 N$7714 "Straight Waveguide" sch_x=111 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3858 N$7715 N$7716 "Straight Waveguide" sch_x=111 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3859 N$7717 N$7718 "Straight Waveguide" sch_x=111 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3860 N$7719 N$7720 "Straight Waveguide" sch_x=111 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3861 N$7721 N$7722 "Straight Waveguide" sch_x=111 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3862 N$7723 N$7724 "Straight Waveguide" sch_x=111 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3863 N$7725 N$7726 "Straight Waveguide" sch_x=111 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3864 N$7727 N$7728 "Straight Waveguide" sch_x=111 sch_y=-23.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3865 N$7729 N$7730 "Straight Waveguide" sch_x=109 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3866 N$7731 N$7732 "Straight Waveguide" sch_x=109 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3867 N$7733 N$7734 "Straight Waveguide" sch_x=109 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3868 N$7735 N$7736 "Straight Waveguide" sch_x=109 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3869 N$7737 N$7738 "Straight Waveguide" sch_x=109 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3870 N$7739 N$7740 "Straight Waveguide" sch_x=109 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3871 N$7741 N$7742 "Straight Waveguide" sch_x=109 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3872 N$7743 N$7744 "Straight Waveguide" sch_x=109 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3873 N$7745 N$7746 "Straight Waveguide" sch_x=109 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3874 N$7747 N$7748 "Straight Waveguide" sch_x=109 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3875 N$7749 N$7750 "Straight Waveguide" sch_x=109 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3876 N$7751 N$7752 "Straight Waveguide" sch_x=109 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3877 N$7753 N$7754 "Straight Waveguide" sch_x=109 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3878 N$7755 N$7756 "Straight Waveguide" sch_x=109 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3879 N$7757 N$7758 "Straight Waveguide" sch_x=109 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3880 N$7759 N$7760 "Straight Waveguide" sch_x=109 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3881 N$7761 N$7762 "Straight Waveguide" sch_x=109 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3882 N$7763 N$7764 "Straight Waveguide" sch_x=109 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3883 N$7765 N$7766 "Straight Waveguide" sch_x=109 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3884 N$7767 N$7768 "Straight Waveguide" sch_x=109 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3885 N$7769 N$7770 "Straight Waveguide" sch_x=109 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3886 N$7771 N$7772 "Straight Waveguide" sch_x=109 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3887 N$7773 N$7774 "Straight Waveguide" sch_x=109 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3888 N$7775 N$7776 "Straight Waveguide" sch_x=109 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3889 N$7777 N$7778 "Straight Waveguide" sch_x=109 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3890 N$7779 N$7780 "Straight Waveguide" sch_x=109 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3891 N$7781 N$7782 "Straight Waveguide" sch_x=109 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3892 N$7783 N$7784 "Straight Waveguide" sch_x=109 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3893 N$7785 N$7786 "Straight Waveguide" sch_x=109 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3894 N$7787 N$7788 "Straight Waveguide" sch_x=109 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3895 N$7789 N$7790 "Straight Waveguide" sch_x=109 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3896 N$7791 N$7792 "Straight Waveguide" sch_x=109 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3897 N$7793 N$7794 "Straight Waveguide" sch_x=109 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3898 N$7795 N$7796 "Straight Waveguide" sch_x=109 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3899 N$7797 N$7798 "Straight Waveguide" sch_x=109 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3900 N$7799 N$7800 "Straight Waveguide" sch_x=109 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3901 N$7801 N$7802 "Straight Waveguide" sch_x=109 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3902 N$7803 N$7804 "Straight Waveguide" sch_x=109 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3903 N$7805 N$7806 "Straight Waveguide" sch_x=109 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3904 N$7807 N$7808 "Straight Waveguide" sch_x=109 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3905 N$7809 N$7810 "Straight Waveguide" sch_x=109 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3906 N$7811 N$7812 "Straight Waveguide" sch_x=109 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3907 N$7813 N$7814 "Straight Waveguide" sch_x=109 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3908 N$7815 N$7816 "Straight Waveguide" sch_x=109 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3909 N$7817 N$7818 "Straight Waveguide" sch_x=109 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3910 N$7819 N$7820 "Straight Waveguide" sch_x=109 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3911 N$7821 N$7822 "Straight Waveguide" sch_x=107 sch_y=21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3912 N$7823 N$7824 "Straight Waveguide" sch_x=107 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3913 N$7825 N$7826 "Straight Waveguide" sch_x=107 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3914 N$7827 N$7828 "Straight Waveguide" sch_x=107 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3915 N$7829 N$7830 "Straight Waveguide" sch_x=107 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3916 N$7831 N$7832 "Straight Waveguide" sch_x=107 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3917 N$7833 N$7834 "Straight Waveguide" sch_x=107 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3918 N$7835 N$7836 "Straight Waveguide" sch_x=107 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3919 N$7837 N$7838 "Straight Waveguide" sch_x=107 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3920 N$7839 N$7840 "Straight Waveguide" sch_x=107 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3921 N$7841 N$7842 "Straight Waveguide" sch_x=107 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3922 N$7843 N$7844 "Straight Waveguide" sch_x=107 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3923 N$7845 N$7846 "Straight Waveguide" sch_x=107 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3924 N$7847 N$7848 "Straight Waveguide" sch_x=107 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3925 N$7849 N$7850 "Straight Waveguide" sch_x=107 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3926 N$7851 N$7852 "Straight Waveguide" sch_x=107 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3927 N$7853 N$7854 "Straight Waveguide" sch_x=107 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3928 N$7855 N$7856 "Straight Waveguide" sch_x=107 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3929 N$7857 N$7858 "Straight Waveguide" sch_x=107 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3930 N$7859 N$7860 "Straight Waveguide" sch_x=107 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3931 N$7861 N$7862 "Straight Waveguide" sch_x=107 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3932 N$7863 N$7864 "Straight Waveguide" sch_x=107 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3933 N$7865 N$7866 "Straight Waveguide" sch_x=107 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3934 N$7867 N$7868 "Straight Waveguide" sch_x=107 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3935 N$7869 N$7870 "Straight Waveguide" sch_x=107 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3936 N$7871 N$7872 "Straight Waveguide" sch_x=107 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3937 N$7873 N$7874 "Straight Waveguide" sch_x=107 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3938 N$7875 N$7876 "Straight Waveguide" sch_x=107 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3939 N$7877 N$7878 "Straight Waveguide" sch_x=107 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3940 N$7879 N$7880 "Straight Waveguide" sch_x=107 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3941 N$7881 N$7882 "Straight Waveguide" sch_x=107 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3942 N$7883 N$7884 "Straight Waveguide" sch_x=107 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3943 N$7885 N$7886 "Straight Waveguide" sch_x=107 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3944 N$7887 N$7888 "Straight Waveguide" sch_x=107 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3945 N$7889 N$7890 "Straight Waveguide" sch_x=107 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3946 N$7891 N$7892 "Straight Waveguide" sch_x=107 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3947 N$7893 N$7894 "Straight Waveguide" sch_x=107 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3948 N$7895 N$7896 "Straight Waveguide" sch_x=107 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3949 N$7897 N$7898 "Straight Waveguide" sch_x=107 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3950 N$7899 N$7900 "Straight Waveguide" sch_x=107 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3951 N$7901 N$7902 "Straight Waveguide" sch_x=107 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3952 N$7903 N$7904 "Straight Waveguide" sch_x=107 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3953 N$7905 N$7906 "Straight Waveguide" sch_x=107 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3954 N$7907 N$7908 "Straight Waveguide" sch_x=107 sch_y=-21.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3955 N$7909 N$7910 "Straight Waveguide" sch_x=105 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3956 N$7911 N$7912 "Straight Waveguide" sch_x=105 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3957 N$7913 N$7914 "Straight Waveguide" sch_x=105 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3958 N$7915 N$7916 "Straight Waveguide" sch_x=105 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3959 N$7917 N$7918 "Straight Waveguide" sch_x=105 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3960 N$7919 N$7920 "Straight Waveguide" sch_x=105 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3961 N$7921 N$7922 "Straight Waveguide" sch_x=105 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3962 N$7923 N$7924 "Straight Waveguide" sch_x=105 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3963 N$7925 N$7926 "Straight Waveguide" sch_x=105 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3964 N$7927 N$7928 "Straight Waveguide" sch_x=105 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3965 N$7929 N$7930 "Straight Waveguide" sch_x=105 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3966 N$7931 N$7932 "Straight Waveguide" sch_x=105 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3967 N$7933 N$7934 "Straight Waveguide" sch_x=105 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3968 N$7935 N$7936 "Straight Waveguide" sch_x=105 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3969 N$7937 N$7938 "Straight Waveguide" sch_x=105 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3970 N$7939 N$7940 "Straight Waveguide" sch_x=105 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3971 N$7941 N$7942 "Straight Waveguide" sch_x=105 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3972 N$7943 N$7944 "Straight Waveguide" sch_x=105 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3973 N$7945 N$7946 "Straight Waveguide" sch_x=105 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3974 N$7947 N$7948 "Straight Waveguide" sch_x=105 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3975 N$7949 N$7950 "Straight Waveguide" sch_x=105 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3976 N$7951 N$7952 "Straight Waveguide" sch_x=105 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3977 N$7953 N$7954 "Straight Waveguide" sch_x=105 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3978 N$7955 N$7956 "Straight Waveguide" sch_x=105 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3979 N$7957 N$7958 "Straight Waveguide" sch_x=105 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3980 N$7959 N$7960 "Straight Waveguide" sch_x=105 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3981 N$7961 N$7962 "Straight Waveguide" sch_x=105 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3982 N$7963 N$7964 "Straight Waveguide" sch_x=105 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3983 N$7965 N$7966 "Straight Waveguide" sch_x=105 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3984 N$7967 N$7968 "Straight Waveguide" sch_x=105 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3985 N$7969 N$7970 "Straight Waveguide" sch_x=105 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3986 N$7971 N$7972 "Straight Waveguide" sch_x=105 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3987 N$7973 N$7974 "Straight Waveguide" sch_x=105 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3988 N$7975 N$7976 "Straight Waveguide" sch_x=105 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3989 N$7977 N$7978 "Straight Waveguide" sch_x=105 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3990 N$7979 N$7980 "Straight Waveguide" sch_x=105 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3991 N$7981 N$7982 "Straight Waveguide" sch_x=105 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3992 N$7983 N$7984 "Straight Waveguide" sch_x=105 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3993 N$7985 N$7986 "Straight Waveguide" sch_x=105 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3994 N$7987 N$7988 "Straight Waveguide" sch_x=105 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3995 N$7989 N$7990 "Straight Waveguide" sch_x=105 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3996 N$7991 N$7992 "Straight Waveguide" sch_x=105 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3997 N$7993 N$7994 "Straight Waveguide" sch_x=103 sch_y=19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3998 N$7995 N$7996 "Straight Waveguide" sch_x=103 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W3999 N$7997 N$7998 "Straight Waveguide" sch_x=103 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4000 N$7999 N$8000 "Straight Waveguide" sch_x=103 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4001 N$8001 N$8002 "Straight Waveguide" sch_x=103 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4002 N$8003 N$8004 "Straight Waveguide" sch_x=103 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4003 N$8005 N$8006 "Straight Waveguide" sch_x=103 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4004 N$8007 N$8008 "Straight Waveguide" sch_x=103 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4005 N$8009 N$8010 "Straight Waveguide" sch_x=103 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4006 N$8011 N$8012 "Straight Waveguide" sch_x=103 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4007 N$8013 N$8014 "Straight Waveguide" sch_x=103 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4008 N$8015 N$8016 "Straight Waveguide" sch_x=103 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4009 N$8017 N$8018 "Straight Waveguide" sch_x=103 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4010 N$8019 N$8020 "Straight Waveguide" sch_x=103 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4011 N$8021 N$8022 "Straight Waveguide" sch_x=103 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4012 N$8023 N$8024 "Straight Waveguide" sch_x=103 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4013 N$8025 N$8026 "Straight Waveguide" sch_x=103 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4014 N$8027 N$8028 "Straight Waveguide" sch_x=103 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4015 N$8029 N$8030 "Straight Waveguide" sch_x=103 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4016 N$8031 N$8032 "Straight Waveguide" sch_x=103 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4017 N$8033 N$8034 "Straight Waveguide" sch_x=103 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4018 N$8035 N$8036 "Straight Waveguide" sch_x=103 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4019 N$8037 N$8038 "Straight Waveguide" sch_x=103 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4020 N$8039 N$8040 "Straight Waveguide" sch_x=103 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4021 N$8041 N$8042 "Straight Waveguide" sch_x=103 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4022 N$8043 N$8044 "Straight Waveguide" sch_x=103 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4023 N$8045 N$8046 "Straight Waveguide" sch_x=103 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4024 N$8047 N$8048 "Straight Waveguide" sch_x=103 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4025 N$8049 N$8050 "Straight Waveguide" sch_x=103 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4026 N$8051 N$8052 "Straight Waveguide" sch_x=103 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4027 N$8053 N$8054 "Straight Waveguide" sch_x=103 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4028 N$8055 N$8056 "Straight Waveguide" sch_x=103 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4029 N$8057 N$8058 "Straight Waveguide" sch_x=103 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4030 N$8059 N$8060 "Straight Waveguide" sch_x=103 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4031 N$8061 N$8062 "Straight Waveguide" sch_x=103 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4032 N$8063 N$8064 "Straight Waveguide" sch_x=103 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4033 N$8065 N$8066 "Straight Waveguide" sch_x=103 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4034 N$8067 N$8068 "Straight Waveguide" sch_x=103 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4035 N$8069 N$8070 "Straight Waveguide" sch_x=103 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4036 N$8071 N$8072 "Straight Waveguide" sch_x=103 sch_y=-19.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4037 N$8073 N$8074 "Straight Waveguide" sch_x=101 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4038 N$8075 N$8076 "Straight Waveguide" sch_x=101 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4039 N$8077 N$8078 "Straight Waveguide" sch_x=101 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4040 N$8079 N$8080 "Straight Waveguide" sch_x=101 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4041 N$8081 N$8082 "Straight Waveguide" sch_x=101 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4042 N$8083 N$8084 "Straight Waveguide" sch_x=101 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4043 N$8085 N$8086 "Straight Waveguide" sch_x=101 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4044 N$8087 N$8088 "Straight Waveguide" sch_x=101 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4045 N$8089 N$8090 "Straight Waveguide" sch_x=101 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4046 N$8091 N$8092 "Straight Waveguide" sch_x=101 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4047 N$8093 N$8094 "Straight Waveguide" sch_x=101 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4048 N$8095 N$8096 "Straight Waveguide" sch_x=101 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4049 N$8097 N$8098 "Straight Waveguide" sch_x=101 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4050 N$8099 N$8100 "Straight Waveguide" sch_x=101 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4051 N$8101 N$8102 "Straight Waveguide" sch_x=101 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4052 N$8103 N$8104 "Straight Waveguide" sch_x=101 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4053 N$8105 N$8106 "Straight Waveguide" sch_x=101 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4054 N$8107 N$8108 "Straight Waveguide" sch_x=101 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4055 N$8109 N$8110 "Straight Waveguide" sch_x=101 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4056 N$8111 N$8112 "Straight Waveguide" sch_x=101 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4057 N$8113 N$8114 "Straight Waveguide" sch_x=101 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4058 N$8115 N$8116 "Straight Waveguide" sch_x=101 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4059 N$8117 N$8118 "Straight Waveguide" sch_x=101 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4060 N$8119 N$8120 "Straight Waveguide" sch_x=101 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4061 N$8121 N$8122 "Straight Waveguide" sch_x=101 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4062 N$8123 N$8124 "Straight Waveguide" sch_x=101 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4063 N$8125 N$8126 "Straight Waveguide" sch_x=101 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4064 N$8127 N$8128 "Straight Waveguide" sch_x=101 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4065 N$8129 N$8130 "Straight Waveguide" sch_x=101 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4066 N$8131 N$8132 "Straight Waveguide" sch_x=101 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4067 N$8133 N$8134 "Straight Waveguide" sch_x=101 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4068 N$8135 N$8136 "Straight Waveguide" sch_x=101 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4069 N$8137 N$8138 "Straight Waveguide" sch_x=101 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4070 N$8139 N$8140 "Straight Waveguide" sch_x=101 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4071 N$8141 N$8142 "Straight Waveguide" sch_x=101 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4072 N$8143 N$8144 "Straight Waveguide" sch_x=101 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4073 N$8145 N$8146 "Straight Waveguide" sch_x=101 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4074 N$8147 N$8148 "Straight Waveguide" sch_x=101 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4075 N$8149 N$8150 "Straight Waveguide" sch_x=99 sch_y=17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4076 N$8151 N$8152 "Straight Waveguide" sch_x=99 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4077 N$8153 N$8154 "Straight Waveguide" sch_x=99 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4078 N$8155 N$8156 "Straight Waveguide" sch_x=99 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4079 N$8157 N$8158 "Straight Waveguide" sch_x=99 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4080 N$8159 N$8160 "Straight Waveguide" sch_x=99 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4081 N$8161 N$8162 "Straight Waveguide" sch_x=99 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4082 N$8163 N$8164 "Straight Waveguide" sch_x=99 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4083 N$8165 N$8166 "Straight Waveguide" sch_x=99 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4084 N$8167 N$8168 "Straight Waveguide" sch_x=99 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4085 N$8169 N$8170 "Straight Waveguide" sch_x=99 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4086 N$8171 N$8172 "Straight Waveguide" sch_x=99 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4087 N$8173 N$8174 "Straight Waveguide" sch_x=99 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4088 N$8175 N$8176 "Straight Waveguide" sch_x=99 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4089 N$8177 N$8178 "Straight Waveguide" sch_x=99 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4090 N$8179 N$8180 "Straight Waveguide" sch_x=99 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4091 N$8181 N$8182 "Straight Waveguide" sch_x=99 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4092 N$8183 N$8184 "Straight Waveguide" sch_x=99 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4093 N$8185 N$8186 "Straight Waveguide" sch_x=99 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4094 N$8187 N$8188 "Straight Waveguide" sch_x=99 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4095 N$8189 N$8190 "Straight Waveguide" sch_x=99 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4096 N$8191 N$8192 "Straight Waveguide" sch_x=99 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4097 N$8193 N$8194 "Straight Waveguide" sch_x=99 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4098 N$8195 N$8196 "Straight Waveguide" sch_x=99 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4099 N$8197 N$8198 "Straight Waveguide" sch_x=99 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4100 N$8199 N$8200 "Straight Waveguide" sch_x=99 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4101 N$8201 N$8202 "Straight Waveguide" sch_x=99 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4102 N$8203 N$8204 "Straight Waveguide" sch_x=99 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4103 N$8205 N$8206 "Straight Waveguide" sch_x=99 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4104 N$8207 N$8208 "Straight Waveguide" sch_x=99 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4105 N$8209 N$8210 "Straight Waveguide" sch_x=99 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4106 N$8211 N$8212 "Straight Waveguide" sch_x=99 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4107 N$8213 N$8214 "Straight Waveguide" sch_x=99 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4108 N$8215 N$8216 "Straight Waveguide" sch_x=99 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4109 N$8217 N$8218 "Straight Waveguide" sch_x=99 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4110 N$8219 N$8220 "Straight Waveguide" sch_x=99 sch_y=-17.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4111 N$8221 N$8222 "Straight Waveguide" sch_x=97 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4112 N$8223 N$8224 "Straight Waveguide" sch_x=97 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4113 N$8225 N$8226 "Straight Waveguide" sch_x=97 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4114 N$8227 N$8228 "Straight Waveguide" sch_x=97 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4115 N$8229 N$8230 "Straight Waveguide" sch_x=97 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4116 N$8231 N$8232 "Straight Waveguide" sch_x=97 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4117 N$8233 N$8234 "Straight Waveguide" sch_x=97 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4118 N$8235 N$8236 "Straight Waveguide" sch_x=97 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4119 N$8237 N$8238 "Straight Waveguide" sch_x=97 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4120 N$8239 N$8240 "Straight Waveguide" sch_x=97 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4121 N$8241 N$8242 "Straight Waveguide" sch_x=97 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4122 N$8243 N$8244 "Straight Waveguide" sch_x=97 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4123 N$8245 N$8246 "Straight Waveguide" sch_x=97 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4124 N$8247 N$8248 "Straight Waveguide" sch_x=97 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4125 N$8249 N$8250 "Straight Waveguide" sch_x=97 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4126 N$8251 N$8252 "Straight Waveguide" sch_x=97 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4127 N$8253 N$8254 "Straight Waveguide" sch_x=97 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4128 N$8255 N$8256 "Straight Waveguide" sch_x=97 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4129 N$8257 N$8258 "Straight Waveguide" sch_x=97 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4130 N$8259 N$8260 "Straight Waveguide" sch_x=97 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4131 N$8261 N$8262 "Straight Waveguide" sch_x=97 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4132 N$8263 N$8264 "Straight Waveguide" sch_x=97 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4133 N$8265 N$8266 "Straight Waveguide" sch_x=97 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4134 N$8267 N$8268 "Straight Waveguide" sch_x=97 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4135 N$8269 N$8270 "Straight Waveguide" sch_x=97 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4136 N$8271 N$8272 "Straight Waveguide" sch_x=97 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4137 N$8273 N$8274 "Straight Waveguide" sch_x=97 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4138 N$8275 N$8276 "Straight Waveguide" sch_x=97 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4139 N$8277 N$8278 "Straight Waveguide" sch_x=97 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4140 N$8279 N$8280 "Straight Waveguide" sch_x=97 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4141 N$8281 N$8282 "Straight Waveguide" sch_x=97 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4142 N$8283 N$8284 "Straight Waveguide" sch_x=97 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4143 N$8285 N$8286 "Straight Waveguide" sch_x=97 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4144 N$8287 N$8288 "Straight Waveguide" sch_x=97 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4145 N$8289 N$8290 "Straight Waveguide" sch_x=95 sch_y=15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4146 N$8291 N$8292 "Straight Waveguide" sch_x=95 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4147 N$8293 N$8294 "Straight Waveguide" sch_x=95 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4148 N$8295 N$8296 "Straight Waveguide" sch_x=95 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4149 N$8297 N$8298 "Straight Waveguide" sch_x=95 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4150 N$8299 N$8300 "Straight Waveguide" sch_x=95 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4151 N$8301 N$8302 "Straight Waveguide" sch_x=95 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4152 N$8303 N$8304 "Straight Waveguide" sch_x=95 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4153 N$8305 N$8306 "Straight Waveguide" sch_x=95 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4154 N$8307 N$8308 "Straight Waveguide" sch_x=95 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4155 N$8309 N$8310 "Straight Waveguide" sch_x=95 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4156 N$8311 N$8312 "Straight Waveguide" sch_x=95 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4157 N$8313 N$8314 "Straight Waveguide" sch_x=95 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4158 N$8315 N$8316 "Straight Waveguide" sch_x=95 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4159 N$8317 N$8318 "Straight Waveguide" sch_x=95 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4160 N$8319 N$8320 "Straight Waveguide" sch_x=95 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4161 N$8321 N$8322 "Straight Waveguide" sch_x=95 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4162 N$8323 N$8324 "Straight Waveguide" sch_x=95 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4163 N$8325 N$8326 "Straight Waveguide" sch_x=95 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4164 N$8327 N$8328 "Straight Waveguide" sch_x=95 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4165 N$8329 N$8330 "Straight Waveguide" sch_x=95 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4166 N$8331 N$8332 "Straight Waveguide" sch_x=95 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4167 N$8333 N$8334 "Straight Waveguide" sch_x=95 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4168 N$8335 N$8336 "Straight Waveguide" sch_x=95 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4169 N$8337 N$8338 "Straight Waveguide" sch_x=95 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4170 N$8339 N$8340 "Straight Waveguide" sch_x=95 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4171 N$8341 N$8342 "Straight Waveguide" sch_x=95 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4172 N$8343 N$8344 "Straight Waveguide" sch_x=95 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4173 N$8345 N$8346 "Straight Waveguide" sch_x=95 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4174 N$8347 N$8348 "Straight Waveguide" sch_x=95 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4175 N$8349 N$8350 "Straight Waveguide" sch_x=95 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4176 N$8351 N$8352 "Straight Waveguide" sch_x=95 sch_y=-15.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4177 N$8353 N$8354 "Straight Waveguide" sch_x=93 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4178 N$8355 N$8356 "Straight Waveguide" sch_x=93 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4179 N$8357 N$8358 "Straight Waveguide" sch_x=93 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4180 N$8359 N$8360 "Straight Waveguide" sch_x=93 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4181 N$8361 N$8362 "Straight Waveguide" sch_x=93 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4182 N$8363 N$8364 "Straight Waveguide" sch_x=93 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4183 N$8365 N$8366 "Straight Waveguide" sch_x=93 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4184 N$8367 N$8368 "Straight Waveguide" sch_x=93 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4185 N$8369 N$8370 "Straight Waveguide" sch_x=93 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4186 N$8371 N$8372 "Straight Waveguide" sch_x=93 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4187 N$8373 N$8374 "Straight Waveguide" sch_x=93 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4188 N$8375 N$8376 "Straight Waveguide" sch_x=93 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4189 N$8377 N$8378 "Straight Waveguide" sch_x=93 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4190 N$8379 N$8380 "Straight Waveguide" sch_x=93 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4191 N$8381 N$8382 "Straight Waveguide" sch_x=93 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4192 N$8383 N$8384 "Straight Waveguide" sch_x=93 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4193 N$8385 N$8386 "Straight Waveguide" sch_x=93 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4194 N$8387 N$8388 "Straight Waveguide" sch_x=93 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4195 N$8389 N$8390 "Straight Waveguide" sch_x=93 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4196 N$8391 N$8392 "Straight Waveguide" sch_x=93 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4197 N$8393 N$8394 "Straight Waveguide" sch_x=93 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4198 N$8395 N$8396 "Straight Waveguide" sch_x=93 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4199 N$8397 N$8398 "Straight Waveguide" sch_x=93 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4200 N$8399 N$8400 "Straight Waveguide" sch_x=93 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4201 N$8401 N$8402 "Straight Waveguide" sch_x=93 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4202 N$8403 N$8404 "Straight Waveguide" sch_x=93 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4203 N$8405 N$8406 "Straight Waveguide" sch_x=93 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4204 N$8407 N$8408 "Straight Waveguide" sch_x=93 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4205 N$8409 N$8410 "Straight Waveguide" sch_x=93 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4206 N$8411 N$8412 "Straight Waveguide" sch_x=93 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4207 N$8413 N$8414 "Straight Waveguide" sch_x=91 sch_y=13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4208 N$8415 N$8416 "Straight Waveguide" sch_x=91 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4209 N$8417 N$8418 "Straight Waveguide" sch_x=91 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4210 N$8419 N$8420 "Straight Waveguide" sch_x=91 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4211 N$8421 N$8422 "Straight Waveguide" sch_x=91 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4212 N$8423 N$8424 "Straight Waveguide" sch_x=91 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4213 N$8425 N$8426 "Straight Waveguide" sch_x=91 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4214 N$8427 N$8428 "Straight Waveguide" sch_x=91 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4215 N$8429 N$8430 "Straight Waveguide" sch_x=91 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4216 N$8431 N$8432 "Straight Waveguide" sch_x=91 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4217 N$8433 N$8434 "Straight Waveguide" sch_x=91 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4218 N$8435 N$8436 "Straight Waveguide" sch_x=91 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4219 N$8437 N$8438 "Straight Waveguide" sch_x=91 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4220 N$8439 N$8440 "Straight Waveguide" sch_x=91 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4221 N$8441 N$8442 "Straight Waveguide" sch_x=91 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4222 N$8443 N$8444 "Straight Waveguide" sch_x=91 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4223 N$8445 N$8446 "Straight Waveguide" sch_x=91 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4224 N$8447 N$8448 "Straight Waveguide" sch_x=91 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4225 N$8449 N$8450 "Straight Waveguide" sch_x=91 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4226 N$8451 N$8452 "Straight Waveguide" sch_x=91 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4227 N$8453 N$8454 "Straight Waveguide" sch_x=91 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4228 N$8455 N$8456 "Straight Waveguide" sch_x=91 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4229 N$8457 N$8458 "Straight Waveguide" sch_x=91 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4230 N$8459 N$8460 "Straight Waveguide" sch_x=91 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4231 N$8461 N$8462 "Straight Waveguide" sch_x=91 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4232 N$8463 N$8464 "Straight Waveguide" sch_x=91 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4233 N$8465 N$8466 "Straight Waveguide" sch_x=91 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4234 N$8467 N$8468 "Straight Waveguide" sch_x=91 sch_y=-13.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4235 N$8469 N$8470 "Straight Waveguide" sch_x=89 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4236 N$8471 N$8472 "Straight Waveguide" sch_x=89 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4237 N$8473 N$8474 "Straight Waveguide" sch_x=89 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4238 N$8475 N$8476 "Straight Waveguide" sch_x=89 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4239 N$8477 N$8478 "Straight Waveguide" sch_x=89 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4240 N$8479 N$8480 "Straight Waveguide" sch_x=89 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4241 N$8481 N$8482 "Straight Waveguide" sch_x=89 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4242 N$8483 N$8484 "Straight Waveguide" sch_x=89 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4243 N$8485 N$8486 "Straight Waveguide" sch_x=89 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4244 N$8487 N$8488 "Straight Waveguide" sch_x=89 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4245 N$8489 N$8490 "Straight Waveguide" sch_x=89 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4246 N$8491 N$8492 "Straight Waveguide" sch_x=89 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4247 N$8493 N$8494 "Straight Waveguide" sch_x=89 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4248 N$8495 N$8496 "Straight Waveguide" sch_x=89 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4249 N$8497 N$8498 "Straight Waveguide" sch_x=89 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4250 N$8499 N$8500 "Straight Waveguide" sch_x=89 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4251 N$8501 N$8502 "Straight Waveguide" sch_x=89 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4252 N$8503 N$8504 "Straight Waveguide" sch_x=89 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4253 N$8505 N$8506 "Straight Waveguide" sch_x=89 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4254 N$8507 N$8508 "Straight Waveguide" sch_x=89 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4255 N$8509 N$8510 "Straight Waveguide" sch_x=89 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4256 N$8511 N$8512 "Straight Waveguide" sch_x=89 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4257 N$8513 N$8514 "Straight Waveguide" sch_x=89 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4258 N$8515 N$8516 "Straight Waveguide" sch_x=89 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4259 N$8517 N$8518 "Straight Waveguide" sch_x=89 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4260 N$8519 N$8520 "Straight Waveguide" sch_x=89 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4261 N$8521 N$8522 "Straight Waveguide" sch_x=87 sch_y=11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4262 N$8523 N$8524 "Straight Waveguide" sch_x=87 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4263 N$8525 N$8526 "Straight Waveguide" sch_x=87 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4264 N$8527 N$8528 "Straight Waveguide" sch_x=87 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4265 N$8529 N$8530 "Straight Waveguide" sch_x=87 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4266 N$8531 N$8532 "Straight Waveguide" sch_x=87 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4267 N$8533 N$8534 "Straight Waveguide" sch_x=87 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4268 N$8535 N$8536 "Straight Waveguide" sch_x=87 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4269 N$8537 N$8538 "Straight Waveguide" sch_x=87 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4270 N$8539 N$8540 "Straight Waveguide" sch_x=87 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4271 N$8541 N$8542 "Straight Waveguide" sch_x=87 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4272 N$8543 N$8544 "Straight Waveguide" sch_x=87 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4273 N$8545 N$8546 "Straight Waveguide" sch_x=87 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4274 N$8547 N$8548 "Straight Waveguide" sch_x=87 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4275 N$8549 N$8550 "Straight Waveguide" sch_x=87 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4276 N$8551 N$8552 "Straight Waveguide" sch_x=87 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4277 N$8553 N$8554 "Straight Waveguide" sch_x=87 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4278 N$8555 N$8556 "Straight Waveguide" sch_x=87 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4279 N$8557 N$8558 "Straight Waveguide" sch_x=87 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4280 N$8559 N$8560 "Straight Waveguide" sch_x=87 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4281 N$8561 N$8562 "Straight Waveguide" sch_x=87 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4282 N$8563 N$8564 "Straight Waveguide" sch_x=87 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4283 N$8565 N$8566 "Straight Waveguide" sch_x=87 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4284 N$8567 N$8568 "Straight Waveguide" sch_x=87 sch_y=-11.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4285 N$8569 N$8570 "Straight Waveguide" sch_x=85 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4286 N$8571 N$8572 "Straight Waveguide" sch_x=85 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4287 N$8573 N$8574 "Straight Waveguide" sch_x=85 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4288 N$8575 N$8576 "Straight Waveguide" sch_x=85 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4289 N$8577 N$8578 "Straight Waveguide" sch_x=85 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4290 N$8579 N$8580 "Straight Waveguide" sch_x=85 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4291 N$8581 N$8582 "Straight Waveguide" sch_x=85 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4292 N$8583 N$8584 "Straight Waveguide" sch_x=85 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4293 N$8585 N$8586 "Straight Waveguide" sch_x=85 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4294 N$8587 N$8588 "Straight Waveguide" sch_x=85 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4295 N$8589 N$8590 "Straight Waveguide" sch_x=85 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4296 N$8591 N$8592 "Straight Waveguide" sch_x=85 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4297 N$8593 N$8594 "Straight Waveguide" sch_x=85 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4298 N$8595 N$8596 "Straight Waveguide" sch_x=85 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4299 N$8597 N$8598 "Straight Waveguide" sch_x=85 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4300 N$8599 N$8600 "Straight Waveguide" sch_x=85 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4301 N$8601 N$8602 "Straight Waveguide" sch_x=85 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4302 N$8603 N$8604 "Straight Waveguide" sch_x=85 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4303 N$8605 N$8606 "Straight Waveguide" sch_x=85 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4304 N$8607 N$8608 "Straight Waveguide" sch_x=85 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4305 N$8609 N$8610 "Straight Waveguide" sch_x=85 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4306 N$8611 N$8612 "Straight Waveguide" sch_x=85 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4307 N$8613 N$8614 "Straight Waveguide" sch_x=83 sch_y=9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4308 N$8615 N$8616 "Straight Waveguide" sch_x=83 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4309 N$8617 N$8618 "Straight Waveguide" sch_x=83 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4310 N$8619 N$8620 "Straight Waveguide" sch_x=83 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4311 N$8621 N$8622 "Straight Waveguide" sch_x=83 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4312 N$8623 N$8624 "Straight Waveguide" sch_x=83 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4313 N$8625 N$8626 "Straight Waveguide" sch_x=83 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4314 N$8627 N$8628 "Straight Waveguide" sch_x=83 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4315 N$8629 N$8630 "Straight Waveguide" sch_x=83 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4316 N$8631 N$8632 "Straight Waveguide" sch_x=83 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4317 N$8633 N$8634 "Straight Waveguide" sch_x=83 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4318 N$8635 N$8636 "Straight Waveguide" sch_x=83 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4319 N$8637 N$8638 "Straight Waveguide" sch_x=83 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4320 N$8639 N$8640 "Straight Waveguide" sch_x=83 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4321 N$8641 N$8642 "Straight Waveguide" sch_x=83 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4322 N$8643 N$8644 "Straight Waveguide" sch_x=83 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4323 N$8645 N$8646 "Straight Waveguide" sch_x=83 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4324 N$8647 N$8648 "Straight Waveguide" sch_x=83 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4325 N$8649 N$8650 "Straight Waveguide" sch_x=83 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4326 N$8651 N$8652 "Straight Waveguide" sch_x=83 sch_y=-9.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4327 N$8653 N$8654 "Straight Waveguide" sch_x=81 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4328 N$8655 N$8656 "Straight Waveguide" sch_x=81 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4329 N$8657 N$8658 "Straight Waveguide" sch_x=81 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4330 N$8659 N$8660 "Straight Waveguide" sch_x=81 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4331 N$8661 N$8662 "Straight Waveguide" sch_x=81 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4332 N$8663 N$8664 "Straight Waveguide" sch_x=81 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4333 N$8665 N$8666 "Straight Waveguide" sch_x=81 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4334 N$8667 N$8668 "Straight Waveguide" sch_x=81 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4335 N$8669 N$8670 "Straight Waveguide" sch_x=81 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4336 N$8671 N$8672 "Straight Waveguide" sch_x=81 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4337 N$8673 N$8674 "Straight Waveguide" sch_x=81 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4338 N$8675 N$8676 "Straight Waveguide" sch_x=81 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4339 N$8677 N$8678 "Straight Waveguide" sch_x=81 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4340 N$8679 N$8680 "Straight Waveguide" sch_x=81 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4341 N$8681 N$8682 "Straight Waveguide" sch_x=81 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4342 N$8683 N$8684 "Straight Waveguide" sch_x=81 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4343 N$8685 N$8686 "Straight Waveguide" sch_x=81 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4344 N$8687 N$8688 "Straight Waveguide" sch_x=81 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4345 N$8689 N$8690 "Straight Waveguide" sch_x=79 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4346 N$8691 N$8692 "Straight Waveguide" sch_x=79 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4347 N$8693 N$8694 "Straight Waveguide" sch_x=79 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4348 N$8695 N$8696 "Straight Waveguide" sch_x=79 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4349 N$8697 N$8698 "Straight Waveguide" sch_x=79 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4350 N$8699 N$8700 "Straight Waveguide" sch_x=79 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4351 N$8701 N$8702 "Straight Waveguide" sch_x=79 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4352 N$8703 N$8704 "Straight Waveguide" sch_x=79 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4353 N$8705 N$8706 "Straight Waveguide" sch_x=79 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4354 N$8707 N$8708 "Straight Waveguide" sch_x=79 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4355 N$8709 N$8710 "Straight Waveguide" sch_x=79 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4356 N$8711 N$8712 "Straight Waveguide" sch_x=79 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4357 N$8713 N$8714 "Straight Waveguide" sch_x=79 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4358 N$8715 N$8716 "Straight Waveguide" sch_x=79 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4359 N$8717 N$8718 "Straight Waveguide" sch_x=79 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4360 N$8719 N$8720 "Straight Waveguide" sch_x=79 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4361 N$8721 N$8722 "Straight Waveguide" sch_x=77 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4362 N$8723 N$8724 "Straight Waveguide" sch_x=77 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4363 N$8725 N$8726 "Straight Waveguide" sch_x=77 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4364 N$8727 N$8728 "Straight Waveguide" sch_x=77 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4365 N$8729 N$8730 "Straight Waveguide" sch_x=77 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4366 N$8731 N$8732 "Straight Waveguide" sch_x=77 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4367 N$8733 N$8734 "Straight Waveguide" sch_x=77 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4368 N$8735 N$8736 "Straight Waveguide" sch_x=77 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4369 N$8737 N$8738 "Straight Waveguide" sch_x=77 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4370 N$8739 N$8740 "Straight Waveguide" sch_x=77 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4371 N$8741 N$8742 "Straight Waveguide" sch_x=77 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4372 N$8743 N$8744 "Straight Waveguide" sch_x=77 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4373 N$8745 N$8746 "Straight Waveguide" sch_x=77 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4374 N$8747 N$8748 "Straight Waveguide" sch_x=77 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4375 N$8749 N$8750 "Straight Waveguide" sch_x=75 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4376 N$8751 N$8752 "Straight Waveguide" sch_x=75 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4377 N$8753 N$8754 "Straight Waveguide" sch_x=75 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4378 N$8755 N$8756 "Straight Waveguide" sch_x=75 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4379 N$8757 N$8758 "Straight Waveguide" sch_x=75 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4380 N$8759 N$8760 "Straight Waveguide" sch_x=75 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4381 N$8761 N$8762 "Straight Waveguide" sch_x=75 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4382 N$8763 N$8764 "Straight Waveguide" sch_x=75 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4383 N$8765 N$8766 "Straight Waveguide" sch_x=75 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4384 N$8767 N$8768 "Straight Waveguide" sch_x=75 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4385 N$8769 N$8770 "Straight Waveguide" sch_x=75 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4386 N$8771 N$8772 "Straight Waveguide" sch_x=75 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4387 N$8773 N$8774 "Straight Waveguide" sch_x=73 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4388 N$8775 N$8776 "Straight Waveguide" sch_x=73 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4389 N$8777 N$8778 "Straight Waveguide" sch_x=73 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4390 N$8779 N$8780 "Straight Waveguide" sch_x=73 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4391 N$8781 N$8782 "Straight Waveguide" sch_x=73 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4392 N$8783 N$8784 "Straight Waveguide" sch_x=73 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4393 N$8785 N$8786 "Straight Waveguide" sch_x=73 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4394 N$8787 N$8788 "Straight Waveguide" sch_x=73 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4395 N$8789 N$8790 "Straight Waveguide" sch_x=73 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4396 N$8791 N$8792 "Straight Waveguide" sch_x=73 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4397 N$8793 N$8794 "Straight Waveguide" sch_x=71 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4398 N$8795 N$8796 "Straight Waveguide" sch_x=71 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4399 N$8797 N$8798 "Straight Waveguide" sch_x=71 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4400 N$8799 N$8800 "Straight Waveguide" sch_x=71 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4401 N$8801 N$8802 "Straight Waveguide" sch_x=71 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4402 N$8803 N$8804 "Straight Waveguide" sch_x=71 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4403 N$8805 N$8806 "Straight Waveguide" sch_x=71 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4404 N$8807 N$8808 "Straight Waveguide" sch_x=71 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4405 N$8809 N$8810 "Straight Waveguide" sch_x=69 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4406 N$8811 N$8812 "Straight Waveguide" sch_x=69 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4407 N$8813 N$8814 "Straight Waveguide" sch_x=69 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4408 N$8815 N$8816 "Straight Waveguide" sch_x=69 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4409 N$8817 N$8818 "Straight Waveguide" sch_x=69 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4410 N$8819 N$8820 "Straight Waveguide" sch_x=69 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4411 N$8821 N$8822 "Straight Waveguide" sch_x=67 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4412 N$8823 N$8824 "Straight Waveguide" sch_x=67 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4413 N$8825 N$8826 "Straight Waveguide" sch_x=67 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4414 N$8827 N$8828 "Straight Waveguide" sch_x=67 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4415 N$8829 N$8830 "Straight Waveguide" sch_x=65 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4416 N$8831 N$8832 "Straight Waveguide" sch_x=65 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4417 N$8834 N$8833 "Straight Waveguide" sch_x=93 sch_y=30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4418 N$8836 N$8835 "Straight Waveguide" sch_x=92 sch_y=29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4419 N$8838 N$8837 "Straight Waveguide" sch_x=91 sch_y=28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4420 N$8840 N$8839 "Straight Waveguide" sch_x=90 sch_y=27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4421 N$8842 N$8841 "Straight Waveguide" sch_x=89 sch_y=26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4422 N$8844 N$8843 "Straight Waveguide" sch_x=88 sch_y=25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4423 N$8846 N$8845 "Straight Waveguide" sch_x=87 sch_y=24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4424 N$8848 N$8847 "Straight Waveguide" sch_x=86 sch_y=23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4425 N$8850 N$8849 "Straight Waveguide" sch_x=85 sch_y=22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4426 N$8852 N$8851 "Straight Waveguide" sch_x=84 sch_y=21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4427 N$8854 N$8853 "Straight Waveguide" sch_x=83 sch_y=20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4428 N$8856 N$8855 "Straight Waveguide" sch_x=82 sch_y=19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4429 N$8858 N$8857 "Straight Waveguide" sch_x=81 sch_y=18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4430 N$8860 N$8859 "Straight Waveguide" sch_x=80 sch_y=17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4431 N$8862 N$8861 "Straight Waveguide" sch_x=79 sch_y=16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4432 N$8864 N$8863 "Straight Waveguide" sch_x=78 sch_y=15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4433 N$8866 N$8865 "Straight Waveguide" sch_x=77 sch_y=14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4434 N$8868 N$8867 "Straight Waveguide" sch_x=76 sch_y=13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4435 N$8870 N$8869 "Straight Waveguide" sch_x=75 sch_y=12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4436 N$8872 N$8871 "Straight Waveguide" sch_x=74 sch_y=11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4437 N$8874 N$8873 "Straight Waveguide" sch_x=73 sch_y=10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4438 N$8876 N$8875 "Straight Waveguide" sch_x=72 sch_y=9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4439 N$8878 N$8877 "Straight Waveguide" sch_x=71 sch_y=8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4440 N$8880 N$8879 "Straight Waveguide" sch_x=70 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4441 N$8882 N$8881 "Straight Waveguide" sch_x=69 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4442 N$8884 N$8883 "Straight Waveguide" sch_x=68 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4443 N$8886 N$8885 "Straight Waveguide" sch_x=67 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4444 N$8888 N$8887 "Straight Waveguide" sch_x=66 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4445 N$8890 N$8889 "Straight Waveguide" sch_x=65 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4446 N$8892 N$8891 "Straight Waveguide" sch_x=64 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4447 N$8894 N$8893 "Straight Waveguide" sch_x=63 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4448 N$8896 N$8895 "Straight Waveguide" sch_x=63 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4449 N$8898 N$8897 "Straight Waveguide" sch_x=64 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4450 N$8900 N$8899 "Straight Waveguide" sch_x=65 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4451 N$8902 N$8901 "Straight Waveguide" sch_x=66 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4452 N$8904 N$8903 "Straight Waveguide" sch_x=67 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4453 N$8906 N$8905 "Straight Waveguide" sch_x=68 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4454 N$8908 N$8907 "Straight Waveguide" sch_x=69 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4455 N$8910 N$8909 "Straight Waveguide" sch_x=70 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4456 N$8912 N$8911 "Straight Waveguide" sch_x=71 sch_y=-8.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4457 N$8914 N$8913 "Straight Waveguide" sch_x=72 sch_y=-9 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4458 N$8916 N$8915 "Straight Waveguide" sch_x=73 sch_y=-10.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4459 N$8918 N$8917 "Straight Waveguide" sch_x=74 sch_y=-11 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4460 N$8920 N$8919 "Straight Waveguide" sch_x=75 sch_y=-12.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4461 N$8922 N$8921 "Straight Waveguide" sch_x=76 sch_y=-13 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4462 N$8924 N$8923 "Straight Waveguide" sch_x=77 sch_y=-14.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4463 N$8926 N$8925 "Straight Waveguide" sch_x=78 sch_y=-15 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4464 N$8928 N$8927 "Straight Waveguide" sch_x=79 sch_y=-16.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4465 N$8930 N$8929 "Straight Waveguide" sch_x=80 sch_y=-17 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4466 N$8932 N$8931 "Straight Waveguide" sch_x=81 sch_y=-18.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4467 N$8934 N$8933 "Straight Waveguide" sch_x=82 sch_y=-19 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4468 N$8936 N$8935 "Straight Waveguide" sch_x=83 sch_y=-20.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4469 N$8938 N$8937 "Straight Waveguide" sch_x=84 sch_y=-21 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4470 N$8940 N$8939 "Straight Waveguide" sch_x=85 sch_y=-22.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4471 N$8942 N$8941 "Straight Waveguide" sch_x=86 sch_y=-23 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4472 N$8944 N$8943 "Straight Waveguide" sch_x=87 sch_y=-24.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4473 N$8946 N$8945 "Straight Waveguide" sch_x=88 sch_y=-25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4474 N$8948 N$8947 "Straight Waveguide" sch_x=89 sch_y=-26.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4475 N$8950 N$8949 "Straight Waveguide" sch_x=90 sch_y=-27 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4476 N$8952 N$8951 "Straight Waveguide" sch_x=91 sch_y=-28.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4477 N$8954 N$8953 "Straight Waveguide" sch_x=92 sch_y=-29 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4478 N$8956 N$8955 "Straight Waveguide" sch_x=93 sch_y=-30.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4479 N$8958 N$8957 "Straight Waveguide" sch_x=94 sch_y=31 sch_r=0 sch_f=false lay_x=0 lay_y=0
   W4480 N$8960 N$8959 "Straight Waveguide" sch_x=94 sch_y=-31 sch_r=0 sch_f=false lay_x=0 lay_y=0
.ends HDBE
* - ONA
.ona input_unit=wavelength input_parameter=center_and_range center=1550e-9
  + range=100e-9 number_of_points=100 
  + minimum_loss=200
  + sensitivity=-200 
  + analysis_type=scattering_data
  + multithreading=user_defined number_of_threads=1 
 + input(1)=HDBE,N$9153
+ input(2)=HDBE,N$9155
+ input(3)=HDBE,N$9157
+ input(4)=HDBE,N$9159
+ input(5)=HDBE,N$9161
+ input(6)=HDBE,N$9163
+ input(7)=HDBE,N$9165
+ input(8)=HDBE,N$9167
+ input(9)=HDBE,N$9169
+ input(10)=HDBE,N$9171
+ input(11)=HDBE,N$9173
+ input(12)=HDBE,N$9175
+ input(13)=HDBE,N$9177
+ input(14)=HDBE,N$9179
+ input(15)=HDBE,N$9181
+ input(16)=HDBE,N$9183
+ input(17)=HDBE,N$9185
+ input(18)=HDBE,N$9187
+ input(19)=HDBE,N$9189
+ input(20)=HDBE,N$9191
+ input(21)=HDBE,N$9193
+ input(22)=HDBE,N$9195
+ input(23)=HDBE,N$9197
+ input(24)=HDBE,N$9199
+ input(25)=HDBE,N$9201
+ input(26)=HDBE,N$9203
+ input(27)=HDBE,N$9205
+ input(28)=HDBE,N$9207
+ input(29)=HDBE,N$9209
+ input(30)=HDBE,N$9211
+ input(31)=HDBE,N$9213
+ input(32)=HDBE,N$9215
  + output=HDBE,N$8961

HDBE  N$8961 N$8963 N$8965 N$8967 N$8969 N$8971 N$8973 N$8975 N$8977 N$8979 N$8981 N$8983 N$8985 N$8987 N$8989 N$8991 N$8993 N$8995 N$8997 N$8999 N$9001 N$9003 N$9005 N$9007 N$9009 N$9011 N$9013 N$9015 N$9017 N$9019 N$9021 N$9023 N$9153 N$9155 N$9157 N$9159 N$9161 N$9163 N$9165 N$9167 N$9169 N$9171 N$9173 N$9175 N$9177 N$9179 N$9181 N$9183 N$9185 N$9187 N$9189 N$9191 N$9193 N$9195 N$9197 N$9199 N$9201 N$9203 N$9205 N$9207 N$9209 N$9211 N$9213 N$9215 HDBE sch_x=0 sch_y=0
*
.end