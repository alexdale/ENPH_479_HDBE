*
* MAIN CELL: Component pathname : root_element
*
   .MODEL MMI_switch_ideal "label 1"="TE" "control"=1
   .MODEL "Waveguide Crossing" "label 1"="TE" "transmission 1"=0.9954054174 "cross talk 1"=0.0001
   + "transmission 2"=1 "cross talk 2"=0 "reflection 1"=0.001
   + "reflection 2"=0 "label 2"="TM" "orthogonal identifier 1"=1
   + "orthogonal identifier 2"=2
   .MODEL "Straight Waveguide" "excess loss temperature sensitivity 2"=0 "label 1"="TE" "orthogonal identifier 1"=1 
   + "loss 1"=0 "number of taps"=64 "dispersion 1"=0 
   + "effective index temperature sensitivity 2"=0 "effective index 2"=1 length=10u 
   + "group index 2"=1 "orthogonal identifier 2"=2 "nominal temperature"=300 
   + "loss 2"=0 "dispersion 2"=0 frequency=193.1T 
   + "digital filter"=0 "run diagnostic"=0 "window function"="rectangular" 
   + "thermal fill factor"=1 "excess loss temperature sensitivity 1"=0 "label 2"="TM" 
   + "thermal effects"=0 "effective index temperature sensitivity 1"=0 "effective index 1"=1 

   S105 N$321 N$322 N$247 N$177 MMI_switch_ideal library="Design kits/capstone" sch_x=-15 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S106 N$323 N$324 N$178 N$179 MMI_switch_ideal library="Design kits/capstone" sch_x=-15 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S107 N$325 N$326 N$180 N$181 MMI_switch_ideal library="Design kits/capstone" sch_x=-15 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S108 N$327 N$328 N$182 N$183 MMI_switch_ideal library="Design kits/capstone" sch_x=-15 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S109 N$329 N$330 N$184 N$185 MMI_switch_ideal library="Design kits/capstone" sch_x=-15 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S110 N$331 N$332 N$186 N$187 MMI_switch_ideal library="Design kits/capstone" sch_x=-15 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S111 N$333 N$334 N$188 N$189 MMI_switch_ideal library="Design kits/capstone" sch_x=-15 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S112 N$335 N$336 N$190 N$248 MMI_switch_ideal library="Design kits/capstone" sch_x=-15 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C113 N$177 N$178 N$233 N$191 "Waveguide Crossing" sch_x=-14 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C114 N$179 N$180 N$192 N$193 "Waveguide Crossing" sch_x=-14 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C115 N$181 N$182 N$194 N$195 "Waveguide Crossing" sch_x=-14 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C116 N$183 N$184 N$196 N$197 "Waveguide Crossing" sch_x=-14 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C117 N$185 N$186 N$198 N$199 "Waveguide Crossing" sch_x=-14 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C118 N$187 N$188 N$200 N$201 "Waveguide Crossing" sch_x=-14 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C119 N$189 N$190 N$202 N$246 "Waveguide Crossing" sch_x=-14 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C120 N$191 N$192 N$234 N$203 "Waveguide Crossing" sch_x=-13 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C121 N$193 N$194 N$204 N$205 "Waveguide Crossing" sch_x=-13 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C122 N$195 N$196 N$206 N$207 "Waveguide Crossing" sch_x=-13 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C123 N$197 N$198 N$208 N$209 "Waveguide Crossing" sch_x=-13 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C124 N$199 N$200 N$210 N$211 "Waveguide Crossing" sch_x=-13 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C125 N$201 N$202 N$212 N$245 "Waveguide Crossing" sch_x=-13 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C126 N$203 N$204 N$235 N$213 "Waveguide Crossing" sch_x=-12 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C127 N$205 N$206 N$214 N$215 "Waveguide Crossing" sch_x=-12 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C128 N$207 N$208 N$216 N$217 "Waveguide Crossing" sch_x=-12 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C129 N$209 N$210 N$218 N$219 "Waveguide Crossing" sch_x=-12 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C130 N$211 N$212 N$220 N$244 "Waveguide Crossing" sch_x=-12 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C131 N$213 N$214 N$236 N$221 "Waveguide Crossing" sch_x=-11 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C132 N$215 N$216 N$222 N$223 "Waveguide Crossing" sch_x=-11 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C133 N$217 N$218 N$224 N$225 "Waveguide Crossing" sch_x=-11 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C134 N$219 N$220 N$226 N$243 "Waveguide Crossing" sch_x=-11 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C135 N$221 N$222 N$237 N$227 "Waveguide Crossing" sch_x=-10 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C136 N$223 N$224 N$228 N$229 "Waveguide Crossing" sch_x=-10 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C137 N$225 N$226 N$230 N$242 "Waveguide Crossing" sch_x=-10 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C138 N$227 N$228 N$238 N$231 "Waveguide Crossing" sch_x=-9 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C139 N$229 N$230 N$232 N$241 "Waveguide Crossing" sch_x=-9 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C140 N$231 N$232 N$239 N$240 "Waveguide Crossing" sch_x=-8 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S85 N$240 N$241 N$155 N$137 MMI_switch_ideal library="Design kits/capstone" sch_x=-7 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S86 N$242 N$243 N$138 N$139 MMI_switch_ideal library="Design kits/capstone" sch_x=-7 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S87 N$244 N$245 N$140 N$141 MMI_switch_ideal library="Design kits/capstone" sch_x=-7 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S88 N$246 N$248 N$142 N$156 MMI_switch_ideal library="Design kits/capstone" sch_x=-7 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C89 N$137 N$138 N$149 N$143 "Waveguide Crossing" sch_x=-6 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C90 N$139 N$140 N$144 N$145 "Waveguide Crossing" sch_x=-6 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C91 N$141 N$142 N$146 N$154 "Waveguide Crossing" sch_x=-6 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C92 N$143 N$144 N$150 N$147 "Waveguide Crossing" sch_x=-5 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C93 N$145 N$146 N$148 N$153 "Waveguide Crossing" sch_x=-5 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C94 N$147 N$148 N$151 N$152 "Waveguide Crossing" sch_x=-4 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S33 N$247 N$233 N$67 N$49 MMI_switch_ideal library="Design kits/capstone" sch_x=-7 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S34 N$234 N$235 N$50 N$51 MMI_switch_ideal library="Design kits/capstone" sch_x=-7 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S35 N$236 N$237 N$52 N$53 MMI_switch_ideal library="Design kits/capstone" sch_x=-7 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S36 N$238 N$239 N$54 N$68 MMI_switch_ideal library="Design kits/capstone" sch_x=-7 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C37 N$49 N$50 N$61 N$55 "Waveguide Crossing" sch_x=-6 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C38 N$51 N$52 N$56 N$57 "Waveguide Crossing" sch_x=-6 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C39 N$53 N$54 N$58 N$66 "Waveguide Crossing" sch_x=-6 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C40 N$55 N$56 N$62 N$59 "Waveguide Crossing" sch_x=-5 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C41 N$57 N$58 N$60 N$65 "Waveguide Crossing" sch_x=-5 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C42 N$59 N$60 N$63 N$64 "Waveguide Crossing" sch_x=-4 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S1 N$67 N$61 N$1 N$2 MMI_switch_ideal library="Design kits/capstone" sch_x=-3 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S2 N$62 N$63 N$3 N$6 MMI_switch_ideal library="Design kits/capstone" sch_x=-3 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S3 N$337 N$1 N$7 N$8 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S4 N$4 N$338 N$9 N$12 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S5 N$339 N$5 N$13 N$14 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S6 N$6 N$340 N$15 N$18 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S7 N$7 N$11 N$19 N$341 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S8 N$10 N$12 N$342 N$20 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S9 N$13 N$17 N$21 N$343 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S10 N$16 N$18 N$344 N$24 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S11 N$19 N$23 N$87 N$81 MMI_switch_ideal library="Design kits/capstone" sch_x=3 sch_y=6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S12 N$22 N$24 N$82 N$83 MMI_switch_ideal library="Design kits/capstone" sch_x=3 sch_y=5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C13 N$2 N$3 N$4 N$5 "Waveguide Crossing" sch_x=-2 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C14 N$8 N$9 N$11 N$10 "Waveguide Crossing" sch_x=0 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C15 N$14 N$15 N$17 N$16 "Waveguide Crossing" sch_x=0 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C16 N$20 N$21 N$23 N$22 "Waveguide Crossing" sch_x=2 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S17 N$64 N$65 N$25 N$26 MMI_switch_ideal library="Design kits/capstone" sch_x=-3 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S18 N$66 N$68 N$27 N$30 MMI_switch_ideal library="Design kits/capstone" sch_x=-3 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S19 N$345 N$25 N$31 N$32 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S20 N$28 N$346 N$33 N$36 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S21 N$347 N$29 N$37 N$38 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S22 N$30 N$348 N$39 N$42 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S23 N$31 N$35 N$43 N$349 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S24 N$34 N$36 N$350 N$44 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S25 N$37 N$41 N$45 N$351 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S26 N$40 N$42 N$352 N$48 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S27 N$43 N$47 N$84 N$85 MMI_switch_ideal library="Design kits/capstone" sch_x=3 sch_y=2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S28 N$46 N$48 N$86 N$88 MMI_switch_ideal library="Design kits/capstone" sch_x=3 sch_y=1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C29 N$26 N$27 N$28 N$29 "Waveguide Crossing" sch_x=-2 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C30 N$32 N$33 N$35 N$34 "Waveguide Crossing" sch_x=0 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C31 N$38 N$39 N$41 N$40 "Waveguide Crossing" sch_x=0 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C32 N$44 N$45 N$47 N$46 "Waveguide Crossing" sch_x=2 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C47 N$81 N$75 N$69 N$70 "Waveguide Crossing" sch_x=6 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C48 N$76 N$77 N$71 N$72 "Waveguide Crossing" sch_x=6 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C49 N$78 N$86 N$73 N$74 "Waveguide Crossing" sch_x=6 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C50 N$82 N$79 N$75 N$76 "Waveguide Crossing" sch_x=5 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C51 N$80 N$85 N$77 N$78 "Waveguide Crossing" sch_x=5 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C52 N$83 N$84 N$79 N$80 "Waveguide Crossing" sch_x=4 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S43 N$87 N$69 N$319 N$305 MMI_switch_ideal library="Design kits/capstone" sch_x=7 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S44 N$70 N$71 N$306 N$307 MMI_switch_ideal library="Design kits/capstone" sch_x=7 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S45 N$72 N$73 N$308 N$309 MMI_switch_ideal library="Design kits/capstone" sch_x=7 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S46 N$74 N$88 N$310 N$311 MMI_switch_ideal library="Design kits/capstone" sch_x=7 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S53 N$155 N$149 N$89 N$90 MMI_switch_ideal library="Design kits/capstone" sch_x=-3 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S54 N$150 N$151 N$91 N$94 MMI_switch_ideal library="Design kits/capstone" sch_x=-3 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S55 N$353 N$89 N$95 N$96 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S56 N$92 N$354 N$97 N$100 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S57 N$355 N$93 N$101 N$102 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S58 N$94 N$356 N$103 N$106 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S59 N$95 N$99 N$107 N$357 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=-0.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S60 N$98 N$100 N$358 N$108 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=-1.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S61 N$101 N$105 N$109 N$359 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=-2.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S62 N$104 N$106 N$360 N$112 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=-3.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S63 N$107 N$111 N$175 N$169 MMI_switch_ideal library="Design kits/capstone" sch_x=3 sch_y=-1.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S64 N$110 N$112 N$170 N$171 MMI_switch_ideal library="Design kits/capstone" sch_x=3 sch_y=-2.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C65 N$90 N$91 N$92 N$93 "Waveguide Crossing" sch_x=-2 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C66 N$96 N$97 N$99 N$98 "Waveguide Crossing" sch_x=0 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C67 N$102 N$103 N$105 N$104 "Waveguide Crossing" sch_x=0 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C68 N$108 N$109 N$111 N$110 "Waveguide Crossing" sch_x=2 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S69 N$152 N$153 N$113 N$114 MMI_switch_ideal library="Design kits/capstone" sch_x=-3 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S70 N$154 N$156 N$115 N$118 MMI_switch_ideal library="Design kits/capstone" sch_x=-3 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S71 N$361 N$113 N$119 N$120 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S72 N$116 N$362 N$121 N$124 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S73 N$363 N$117 N$125 N$126 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S74 N$118 N$364 N$127 N$130 MMI_switch_ideal library="Design kits/capstone" sch_x=-1 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S75 N$119 N$123 N$131 N$365 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=-4.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S76 N$122 N$124 N$366 N$132 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=-5.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S77 N$125 N$129 N$133 N$367 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=-6.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S78 N$128 N$130 N$368 N$136 MMI_switch_ideal library="Design kits/capstone" sch_x=1 sch_y=-7.5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S79 N$131 N$135 N$172 N$173 MMI_switch_ideal library="Design kits/capstone" sch_x=3 sch_y=-5.25 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S80 N$134 N$136 N$174 N$176 MMI_switch_ideal library="Design kits/capstone" sch_x=3 sch_y=-6.75 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C81 N$114 N$115 N$116 N$117 "Waveguide Crossing" sch_x=-2 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C82 N$120 N$121 N$123 N$122 "Waveguide Crossing" sch_x=0 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C83 N$126 N$127 N$129 N$128 "Waveguide Crossing" sch_x=0 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C84 N$132 N$133 N$135 N$134 "Waveguide Crossing" sch_x=2 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C99 N$169 N$163 N$157 N$158 "Waveguide Crossing" sch_x=6 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C100 N$164 N$165 N$159 N$160 "Waveguide Crossing" sch_x=6 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C101 N$166 N$174 N$161 N$162 "Waveguide Crossing" sch_x=6 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C102 N$170 N$167 N$163 N$164 "Waveguide Crossing" sch_x=5 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C103 N$168 N$173 N$165 N$166 "Waveguide Crossing" sch_x=5 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C104 N$171 N$172 N$167 N$168 "Waveguide Crossing" sch_x=4 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S95 N$175 N$157 N$312 N$313 MMI_switch_ideal library="Design kits/capstone" sch_x=7 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S96 N$158 N$159 N$314 N$315 MMI_switch_ideal library="Design kits/capstone" sch_x=7 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S97 N$160 N$161 N$316 N$317 MMI_switch_ideal library="Design kits/capstone" sch_x=7 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S98 N$162 N$176 N$318 N$320 MMI_switch_ideal library="Design kits/capstone" sch_x=7 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C149 N$305 N$263 N$249 N$250 "Waveguide Crossing" sch_x=14 sch_y=6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C150 N$264 N$265 N$251 N$252 "Waveguide Crossing" sch_x=14 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C151 N$266 N$267 N$253 N$254 "Waveguide Crossing" sch_x=14 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C152 N$268 N$269 N$255 N$256 "Waveguide Crossing" sch_x=14 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C153 N$270 N$271 N$257 N$258 "Waveguide Crossing" sch_x=14 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C154 N$272 N$273 N$259 N$260 "Waveguide Crossing" sch_x=14 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C155 N$274 N$318 N$261 N$262 "Waveguide Crossing" sch_x=14 sch_y=-6 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C156 N$306 N$275 N$263 N$264 "Waveguide Crossing" sch_x=13 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C157 N$276 N$277 N$265 N$266 "Waveguide Crossing" sch_x=13 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C158 N$278 N$279 N$267 N$268 "Waveguide Crossing" sch_x=13 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C159 N$280 N$281 N$269 N$270 "Waveguide Crossing" sch_x=13 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C160 N$282 N$283 N$271 N$272 "Waveguide Crossing" sch_x=13 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C161 N$284 N$317 N$273 N$274 "Waveguide Crossing" sch_x=13 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C162 N$307 N$285 N$275 N$276 "Waveguide Crossing" sch_x=12 sch_y=4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C163 N$286 N$287 N$277 N$278 "Waveguide Crossing" sch_x=12 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C164 N$288 N$289 N$279 N$280 "Waveguide Crossing" sch_x=12 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C165 N$290 N$291 N$281 N$282 "Waveguide Crossing" sch_x=12 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C166 N$292 N$316 N$283 N$284 "Waveguide Crossing" sch_x=12 sch_y=-4 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C167 N$308 N$293 N$285 N$286 "Waveguide Crossing" sch_x=11 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C168 N$294 N$295 N$287 N$288 "Waveguide Crossing" sch_x=11 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C169 N$296 N$297 N$289 N$290 "Waveguide Crossing" sch_x=11 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C170 N$298 N$315 N$291 N$292 "Waveguide Crossing" sch_x=11 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C171 N$309 N$299 N$293 N$294 "Waveguide Crossing" sch_x=10 sch_y=2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C172 N$300 N$301 N$295 N$296 "Waveguide Crossing" sch_x=10 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C173 N$302 N$314 N$297 N$298 "Waveguide Crossing" sch_x=10 sch_y=-2 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C174 N$310 N$303 N$299 N$300 "Waveguide Crossing" sch_x=9 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C175 N$304 N$313 N$301 N$302 "Waveguide Crossing" sch_x=9 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   C176 N$311 N$312 N$303 N$304 "Waveguide Crossing" sch_x=8 sch_y=0 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S141 N$319 N$249 N$369 N$370 MMI_switch_ideal library="Design kits/capstone" sch_x=15 sch_y=7 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S142 N$250 N$251 N$371 N$372 MMI_switch_ideal library="Design kits/capstone" sch_x=15 sch_y=5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S143 N$252 N$253 N$373 N$374 MMI_switch_ideal library="Design kits/capstone" sch_x=15 sch_y=3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S144 N$254 N$255 N$375 N$376 MMI_switch_ideal library="Design kits/capstone" sch_x=15 sch_y=1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S145 N$256 N$257 N$377 N$378 MMI_switch_ideal library="Design kits/capstone" sch_x=15 sch_y=-1 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S146 N$258 N$259 N$379 N$380 MMI_switch_ideal library="Design kits/capstone" sch_x=15 sch_y=-3 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S147 N$260 N$261 N$381 N$382 MMI_switch_ideal library="Design kits/capstone" sch_x=15 sch_y=-5 sch_r=0 sch_f=false lay_x=0 lay_y=0
   S148 N$262 N$320 N$383 N$384 MMI_switch_ideal library="Design kits/capstone" sch_x=15 sch_y=-7 sch_r=0 sch_f=false lay_x=0 lay_y=0
